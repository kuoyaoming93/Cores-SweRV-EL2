module ffinv_lut3 #(
) (
    input [31:0]          inv_in,             // Entrada 1
    output [31:0]         out                 // Salida normal
);

    reg [11:0] mem [0:4095];

    assign out = {20'b0,mem[inv_in[11:0]]};

    assign mem[0] = 12'd4095;
    assign mem[1] = 12'd4094;
    assign mem[2] = 12'd4093;
    assign mem[3] = 12'd4092;
    assign mem[4] = 12'd4091;
    assign mem[5] = 12'd4090;
    assign mem[6] = 12'd4089;
    assign mem[7] = 12'd4088;
    assign mem[8] = 12'd4087;
    assign mem[9] = 12'd4086;
    assign mem[10] = 12'd4085;
    assign mem[11] = 12'd4084;
    assign mem[12] = 12'd4083;
    assign mem[13] = 12'd4082;
    assign mem[14] = 12'd4081;
    assign mem[15] = 12'd4080;
    assign mem[16] = 12'd4079;
    assign mem[17] = 12'd4078;
    assign mem[18] = 12'd4077;
    assign mem[19] = 12'd4076;
    assign mem[20] = 12'd4075;
    assign mem[21] = 12'd4074;
    assign mem[22] = 12'd4073;
    assign mem[23] = 12'd4072;
    assign mem[24] = 12'd4071;
    assign mem[25] = 12'd4070;
    assign mem[26] = 12'd4069;
    assign mem[27] = 12'd4068;
    assign mem[28] = 12'd4067;
    assign mem[29] = 12'd4066;
    assign mem[30] = 12'd4065;
    assign mem[31] = 12'd4064;
    assign mem[32] = 12'd4063;
    assign mem[33] = 12'd4062;
    assign mem[34] = 12'd4061;
    assign mem[35] = 12'd4060;
    assign mem[36] = 12'd4059;
    assign mem[37] = 12'd4058;
    assign mem[38] = 12'd4057;
    assign mem[39] = 12'd4056;
    assign mem[40] = 12'd4055;
    assign mem[41] = 12'd4054;
    assign mem[42] = 12'd4053;
    assign mem[43] = 12'd4052;
    assign mem[44] = 12'd4051;
    assign mem[45] = 12'd4050;
    assign mem[46] = 12'd4049;
    assign mem[47] = 12'd4048;
    assign mem[48] = 12'd4047;
    assign mem[49] = 12'd4046;
    assign mem[50] = 12'd4045;
    assign mem[51] = 12'd4044;
    assign mem[52] = 12'd4043;
    assign mem[53] = 12'd4042;
    assign mem[54] = 12'd4041;
    assign mem[55] = 12'd4040;
    assign mem[56] = 12'd4039;
    assign mem[57] = 12'd4038;
    assign mem[58] = 12'd4037;
    assign mem[59] = 12'd4036;
    assign mem[60] = 12'd4035;
    assign mem[61] = 12'd4034;
    assign mem[62] = 12'd4033;
    assign mem[63] = 12'd4032;
    assign mem[64] = 12'd4031;
    assign mem[65] = 12'd4030;
    assign mem[66] = 12'd4029;
    assign mem[67] = 12'd4028;
    assign mem[68] = 12'd4027;
    assign mem[69] = 12'd4026;
    assign mem[70] = 12'd4025;
    assign mem[71] = 12'd4024;
    assign mem[72] = 12'd4023;
    assign mem[73] = 12'd4022;
    assign mem[74] = 12'd4021;
    assign mem[75] = 12'd4020;
    assign mem[76] = 12'd4019;
    assign mem[77] = 12'd4018;
    assign mem[78] = 12'd4017;
    assign mem[79] = 12'd4016;
    assign mem[80] = 12'd4015;
    assign mem[81] = 12'd4014;
    assign mem[82] = 12'd4013;
    assign mem[83] = 12'd4012;
    assign mem[84] = 12'd4011;
    assign mem[85] = 12'd4010;
    assign mem[86] = 12'd4009;
    assign mem[87] = 12'd4008;
    assign mem[88] = 12'd4007;
    assign mem[89] = 12'd4006;
    assign mem[90] = 12'd4005;
    assign mem[91] = 12'd4004;
    assign mem[92] = 12'd4003;
    assign mem[93] = 12'd4002;
    assign mem[94] = 12'd4001;
    assign mem[95] = 12'd4000;
    assign mem[96] = 12'd3999;
    assign mem[97] = 12'd3998;
    assign mem[98] = 12'd3997;
    assign mem[99] = 12'd3996;
    assign mem[100] = 12'd3995;
    assign mem[101] = 12'd3994;
    assign mem[102] = 12'd3993;
    assign mem[103] = 12'd3992;
    assign mem[104] = 12'd3991;
    assign mem[105] = 12'd3990;
    assign mem[106] = 12'd3989;
    assign mem[107] = 12'd3988;
    assign mem[108] = 12'd3987;
    assign mem[109] = 12'd3986;
    assign mem[110] = 12'd3985;
    assign mem[111] = 12'd3984;
    assign mem[112] = 12'd3983;
    assign mem[113] = 12'd3982;
    assign mem[114] = 12'd3981;
    assign mem[115] = 12'd3980;
    assign mem[116] = 12'd3979;
    assign mem[117] = 12'd3978;
    assign mem[118] = 12'd3977;
    assign mem[119] = 12'd3976;
    assign mem[120] = 12'd3975;
    assign mem[121] = 12'd3974;
    assign mem[122] = 12'd3973;
    assign mem[123] = 12'd3972;
    assign mem[124] = 12'd3971;
    assign mem[125] = 12'd3970;
    assign mem[126] = 12'd3969;
    assign mem[127] = 12'd3968;
    assign mem[128] = 12'd3967;
    assign mem[129] = 12'd3966;
    assign mem[130] = 12'd3965;
    assign mem[131] = 12'd3964;
    assign mem[132] = 12'd3963;
    assign mem[133] = 12'd3962;
    assign mem[134] = 12'd3961;
    assign mem[135] = 12'd3960;
    assign mem[136] = 12'd3959;
    assign mem[137] = 12'd3958;
    assign mem[138] = 12'd3957;
    assign mem[139] = 12'd3956;
    assign mem[140] = 12'd3955;
    assign mem[141] = 12'd3954;
    assign mem[142] = 12'd3953;
    assign mem[143] = 12'd3952;
    assign mem[144] = 12'd3951;
    assign mem[145] = 12'd3950;
    assign mem[146] = 12'd3949;
    assign mem[147] = 12'd3948;
    assign mem[148] = 12'd3947;
    assign mem[149] = 12'd3946;
    assign mem[150] = 12'd3945;
    assign mem[151] = 12'd3944;
    assign mem[152] = 12'd3943;
    assign mem[153] = 12'd3942;
    assign mem[154] = 12'd3941;
    assign mem[155] = 12'd3940;
    assign mem[156] = 12'd3939;
    assign mem[157] = 12'd3938;
    assign mem[158] = 12'd3937;
    assign mem[159] = 12'd3936;
    assign mem[160] = 12'd3935;
    assign mem[161] = 12'd3934;
    assign mem[162] = 12'd3933;
    assign mem[163] = 12'd3932;
    assign mem[164] = 12'd3931;
    assign mem[165] = 12'd3930;
    assign mem[166] = 12'd3929;
    assign mem[167] = 12'd3928;
    assign mem[168] = 12'd3927;
    assign mem[169] = 12'd3926;
    assign mem[170] = 12'd3925;
    assign mem[171] = 12'd3924;
    assign mem[172] = 12'd3923;
    assign mem[173] = 12'd3922;
    assign mem[174] = 12'd3921;
    assign mem[175] = 12'd3920;
    assign mem[176] = 12'd3919;
    assign mem[177] = 12'd3918;
    assign mem[178] = 12'd3917;
    assign mem[179] = 12'd3916;
    assign mem[180] = 12'd3915;
    assign mem[181] = 12'd3914;
    assign mem[182] = 12'd3913;
    assign mem[183] = 12'd3912;
    assign mem[184] = 12'd3911;
    assign mem[185] = 12'd3910;
    assign mem[186] = 12'd3909;
    assign mem[187] = 12'd3908;
    assign mem[188] = 12'd3907;
    assign mem[189] = 12'd3906;
    assign mem[190] = 12'd3905;
    assign mem[191] = 12'd3904;
    assign mem[192] = 12'd3903;
    assign mem[193] = 12'd3902;
    assign mem[194] = 12'd3901;
    assign mem[195] = 12'd3900;
    assign mem[196] = 12'd3899;
    assign mem[197] = 12'd3898;
    assign mem[198] = 12'd3897;
    assign mem[199] = 12'd3896;
    assign mem[200] = 12'd3895;
    assign mem[201] = 12'd3894;
    assign mem[202] = 12'd3893;
    assign mem[203] = 12'd3892;
    assign mem[204] = 12'd3891;
    assign mem[205] = 12'd3890;
    assign mem[206] = 12'd3889;
    assign mem[207] = 12'd3888;
    assign mem[208] = 12'd3887;
    assign mem[209] = 12'd3886;
    assign mem[210] = 12'd3885;
    assign mem[211] = 12'd3884;
    assign mem[212] = 12'd3883;
    assign mem[213] = 12'd3882;
    assign mem[214] = 12'd3881;
    assign mem[215] = 12'd3880;
    assign mem[216] = 12'd3879;
    assign mem[217] = 12'd3878;
    assign mem[218] = 12'd3877;
    assign mem[219] = 12'd3876;
    assign mem[220] = 12'd3875;
    assign mem[221] = 12'd3874;
    assign mem[222] = 12'd3873;
    assign mem[223] = 12'd3872;
    assign mem[224] = 12'd3871;
    assign mem[225] = 12'd3870;
    assign mem[226] = 12'd3869;
    assign mem[227] = 12'd3868;
    assign mem[228] = 12'd3867;
    assign mem[229] = 12'd3866;
    assign mem[230] = 12'd3865;
    assign mem[231] = 12'd3864;
    assign mem[232] = 12'd3863;
    assign mem[233] = 12'd3862;
    assign mem[234] = 12'd3861;
    assign mem[235] = 12'd3860;
    assign mem[236] = 12'd3859;
    assign mem[237] = 12'd3858;
    assign mem[238] = 12'd3857;
    assign mem[239] = 12'd3856;
    assign mem[240] = 12'd3855;
    assign mem[241] = 12'd3854;
    assign mem[242] = 12'd3853;
    assign mem[243] = 12'd3852;
    assign mem[244] = 12'd3851;
    assign mem[245] = 12'd3850;
    assign mem[246] = 12'd3849;
    assign mem[247] = 12'd3848;
    assign mem[248] = 12'd3847;
    assign mem[249] = 12'd3846;
    assign mem[250] = 12'd3845;
    assign mem[251] = 12'd3844;
    assign mem[252] = 12'd3843;
    assign mem[253] = 12'd3842;
    assign mem[254] = 12'd3841;
    assign mem[255] = 12'd3840;
    assign mem[256] = 12'd3839;
    assign mem[257] = 12'd3838;
    assign mem[258] = 12'd3837;
    assign mem[259] = 12'd3836;
    assign mem[260] = 12'd3835;
    assign mem[261] = 12'd3834;
    assign mem[262] = 12'd3833;
    assign mem[263] = 12'd3832;
    assign mem[264] = 12'd3831;
    assign mem[265] = 12'd3830;
    assign mem[266] = 12'd3829;
    assign mem[267] = 12'd3828;
    assign mem[268] = 12'd3827;
    assign mem[269] = 12'd3826;
    assign mem[270] = 12'd3825;
    assign mem[271] = 12'd3824;
    assign mem[272] = 12'd3823;
    assign mem[273] = 12'd3822;
    assign mem[274] = 12'd3821;
    assign mem[275] = 12'd3820;
    assign mem[276] = 12'd3819;
    assign mem[277] = 12'd3818;
    assign mem[278] = 12'd3817;
    assign mem[279] = 12'd3816;
    assign mem[280] = 12'd3815;
    assign mem[281] = 12'd3814;
    assign mem[282] = 12'd3813;
    assign mem[283] = 12'd3812;
    assign mem[284] = 12'd3811;
    assign mem[285] = 12'd3810;
    assign mem[286] = 12'd3809;
    assign mem[287] = 12'd3808;
    assign mem[288] = 12'd3807;
    assign mem[289] = 12'd3806;
    assign mem[290] = 12'd3805;
    assign mem[291] = 12'd3804;
    assign mem[292] = 12'd3803;
    assign mem[293] = 12'd3802;
    assign mem[294] = 12'd3801;
    assign mem[295] = 12'd3800;
    assign mem[296] = 12'd3799;
    assign mem[297] = 12'd3798;
    assign mem[298] = 12'd3797;
    assign mem[299] = 12'd3796;
    assign mem[300] = 12'd3795;
    assign mem[301] = 12'd3794;
    assign mem[302] = 12'd3793;
    assign mem[303] = 12'd3792;
    assign mem[304] = 12'd3791;
    assign mem[305] = 12'd3790;
    assign mem[306] = 12'd3789;
    assign mem[307] = 12'd3788;
    assign mem[308] = 12'd3787;
    assign mem[309] = 12'd3786;
    assign mem[310] = 12'd3785;
    assign mem[311] = 12'd3784;
    assign mem[312] = 12'd3783;
    assign mem[313] = 12'd3782;
    assign mem[314] = 12'd3781;
    assign mem[315] = 12'd3780;
    assign mem[316] = 12'd3779;
    assign mem[317] = 12'd3778;
    assign mem[318] = 12'd3777;
    assign mem[319] = 12'd3776;
    assign mem[320] = 12'd3775;
    assign mem[321] = 12'd3774;
    assign mem[322] = 12'd3773;
    assign mem[323] = 12'd3772;
    assign mem[324] = 12'd3771;
    assign mem[325] = 12'd3770;
    assign mem[326] = 12'd3769;
    assign mem[327] = 12'd3768;
    assign mem[328] = 12'd3767;
    assign mem[329] = 12'd3766;
    assign mem[330] = 12'd3765;
    assign mem[331] = 12'd3764;
    assign mem[332] = 12'd3763;
    assign mem[333] = 12'd3762;
    assign mem[334] = 12'd3761;
    assign mem[335] = 12'd3760;
    assign mem[336] = 12'd3759;
    assign mem[337] = 12'd3758;
    assign mem[338] = 12'd3757;
    assign mem[339] = 12'd3756;
    assign mem[340] = 12'd3755;
    assign mem[341] = 12'd3754;
    assign mem[342] = 12'd3753;
    assign mem[343] = 12'd3752;
    assign mem[344] = 12'd3751;
    assign mem[345] = 12'd3750;
    assign mem[346] = 12'd3749;
    assign mem[347] = 12'd3748;
    assign mem[348] = 12'd3747;
    assign mem[349] = 12'd3746;
    assign mem[350] = 12'd3745;
    assign mem[351] = 12'd3744;
    assign mem[352] = 12'd3743;
    assign mem[353] = 12'd3742;
    assign mem[354] = 12'd3741;
    assign mem[355] = 12'd3740;
    assign mem[356] = 12'd3739;
    assign mem[357] = 12'd3738;
    assign mem[358] = 12'd3737;
    assign mem[359] = 12'd3736;
    assign mem[360] = 12'd3735;
    assign mem[361] = 12'd3734;
    assign mem[362] = 12'd3733;
    assign mem[363] = 12'd3732;
    assign mem[364] = 12'd3731;
    assign mem[365] = 12'd3730;
    assign mem[366] = 12'd3729;
    assign mem[367] = 12'd3728;
    assign mem[368] = 12'd3727;
    assign mem[369] = 12'd3726;
    assign mem[370] = 12'd3725;
    assign mem[371] = 12'd3724;
    assign mem[372] = 12'd3723;
    assign mem[373] = 12'd3722;
    assign mem[374] = 12'd3721;
    assign mem[375] = 12'd3720;
    assign mem[376] = 12'd3719;
    assign mem[377] = 12'd3718;
    assign mem[378] = 12'd3717;
    assign mem[379] = 12'd3716;
    assign mem[380] = 12'd3715;
    assign mem[381] = 12'd3714;
    assign mem[382] = 12'd3713;
    assign mem[383] = 12'd3712;
    assign mem[384] = 12'd3711;
    assign mem[385] = 12'd3710;
    assign mem[386] = 12'd3709;
    assign mem[387] = 12'd3708;
    assign mem[388] = 12'd3707;
    assign mem[389] = 12'd3706;
    assign mem[390] = 12'd3705;
    assign mem[391] = 12'd3704;
    assign mem[392] = 12'd3703;
    assign mem[393] = 12'd3702;
    assign mem[394] = 12'd3701;
    assign mem[395] = 12'd3700;
    assign mem[396] = 12'd3699;
    assign mem[397] = 12'd3698;
    assign mem[398] = 12'd3697;
    assign mem[399] = 12'd3696;
    assign mem[400] = 12'd3695;
    assign mem[401] = 12'd3694;
    assign mem[402] = 12'd3693;
    assign mem[403] = 12'd3692;
    assign mem[404] = 12'd3691;
    assign mem[405] = 12'd3690;
    assign mem[406] = 12'd3689;
    assign mem[407] = 12'd3688;
    assign mem[408] = 12'd3687;
    assign mem[409] = 12'd3686;
    assign mem[410] = 12'd3685;
    assign mem[411] = 12'd3684;
    assign mem[412] = 12'd3683;
    assign mem[413] = 12'd3682;
    assign mem[414] = 12'd3681;
    assign mem[415] = 12'd3680;
    assign mem[416] = 12'd3679;
    assign mem[417] = 12'd3678;
    assign mem[418] = 12'd3677;
    assign mem[419] = 12'd3676;
    assign mem[420] = 12'd3675;
    assign mem[421] = 12'd3674;
    assign mem[422] = 12'd3673;
    assign mem[423] = 12'd3672;
    assign mem[424] = 12'd3671;
    assign mem[425] = 12'd3670;
    assign mem[426] = 12'd3669;
    assign mem[427] = 12'd3668;
    assign mem[428] = 12'd3667;
    assign mem[429] = 12'd3666;
    assign mem[430] = 12'd3665;
    assign mem[431] = 12'd3664;
    assign mem[432] = 12'd3663;
    assign mem[433] = 12'd3662;
    assign mem[434] = 12'd3661;
    assign mem[435] = 12'd3660;
    assign mem[436] = 12'd3659;
    assign mem[437] = 12'd3658;
    assign mem[438] = 12'd3657;
    assign mem[439] = 12'd3656;
    assign mem[440] = 12'd3655;
    assign mem[441] = 12'd3654;
    assign mem[442] = 12'd3653;
    assign mem[443] = 12'd3652;
    assign mem[444] = 12'd3651;
    assign mem[445] = 12'd3650;
    assign mem[446] = 12'd3649;
    assign mem[447] = 12'd3648;
    assign mem[448] = 12'd3647;
    assign mem[449] = 12'd3646;
    assign mem[450] = 12'd3645;
    assign mem[451] = 12'd3644;
    assign mem[452] = 12'd3643;
    assign mem[453] = 12'd3642;
    assign mem[454] = 12'd3641;
    assign mem[455] = 12'd3640;
    assign mem[456] = 12'd3639;
    assign mem[457] = 12'd3638;
    assign mem[458] = 12'd3637;
    assign mem[459] = 12'd3636;
    assign mem[460] = 12'd3635;
    assign mem[461] = 12'd3634;
    assign mem[462] = 12'd3633;
    assign mem[463] = 12'd3632;
    assign mem[464] = 12'd3631;
    assign mem[465] = 12'd3630;
    assign mem[466] = 12'd3629;
    assign mem[467] = 12'd3628;
    assign mem[468] = 12'd3627;
    assign mem[469] = 12'd3626;
    assign mem[470] = 12'd3625;
    assign mem[471] = 12'd3624;
    assign mem[472] = 12'd3623;
    assign mem[473] = 12'd3622;
    assign mem[474] = 12'd3621;
    assign mem[475] = 12'd3620;
    assign mem[476] = 12'd3619;
    assign mem[477] = 12'd3618;
    assign mem[478] = 12'd3617;
    assign mem[479] = 12'd3616;
    assign mem[480] = 12'd3615;
    assign mem[481] = 12'd3614;
    assign mem[482] = 12'd3613;
    assign mem[483] = 12'd3612;
    assign mem[484] = 12'd3611;
    assign mem[485] = 12'd3610;
    assign mem[486] = 12'd3609;
    assign mem[487] = 12'd3608;
    assign mem[488] = 12'd3607;
    assign mem[489] = 12'd3606;
    assign mem[490] = 12'd3605;
    assign mem[491] = 12'd3604;
    assign mem[492] = 12'd3603;
    assign mem[493] = 12'd3602;
    assign mem[494] = 12'd3601;
    assign mem[495] = 12'd3600;
    assign mem[496] = 12'd3599;
    assign mem[497] = 12'd3598;
    assign mem[498] = 12'd3597;
    assign mem[499] = 12'd3596;
    assign mem[500] = 12'd3595;
    assign mem[501] = 12'd3594;
    assign mem[502] = 12'd3593;
    assign mem[503] = 12'd3592;
    assign mem[504] = 12'd3591;
    assign mem[505] = 12'd3590;
    assign mem[506] = 12'd3589;
    assign mem[507] = 12'd3588;
    assign mem[508] = 12'd3587;
    assign mem[509] = 12'd3586;
    assign mem[510] = 12'd3585;
    assign mem[511] = 12'd3584;
    assign mem[512] = 12'd3583;
    assign mem[513] = 12'd3582;
    assign mem[514] = 12'd3581;
    assign mem[515] = 12'd3580;
    assign mem[516] = 12'd3579;
    assign mem[517] = 12'd3578;
    assign mem[518] = 12'd3577;
    assign mem[519] = 12'd3576;
    assign mem[520] = 12'd3575;
    assign mem[521] = 12'd3574;
    assign mem[522] = 12'd3573;
    assign mem[523] = 12'd3572;
    assign mem[524] = 12'd3571;
    assign mem[525] = 12'd3570;
    assign mem[526] = 12'd3569;
    assign mem[527] = 12'd3568;
    assign mem[528] = 12'd3567;
    assign mem[529] = 12'd3566;
    assign mem[530] = 12'd3565;
    assign mem[531] = 12'd3564;
    assign mem[532] = 12'd3563;
    assign mem[533] = 12'd3562;
    assign mem[534] = 12'd3561;
    assign mem[535] = 12'd3560;
    assign mem[536] = 12'd3559;
    assign mem[537] = 12'd3558;
    assign mem[538] = 12'd3557;
    assign mem[539] = 12'd3556;
    assign mem[540] = 12'd3555;
    assign mem[541] = 12'd3554;
    assign mem[542] = 12'd3553;
    assign mem[543] = 12'd3552;
    assign mem[544] = 12'd3551;
    assign mem[545] = 12'd3550;
    assign mem[546] = 12'd3549;
    assign mem[547] = 12'd3548;
    assign mem[548] = 12'd3547;
    assign mem[549] = 12'd3546;
    assign mem[550] = 12'd3545;
    assign mem[551] = 12'd3544;
    assign mem[552] = 12'd3543;
    assign mem[553] = 12'd3542;
    assign mem[554] = 12'd3541;
    assign mem[555] = 12'd3540;
    assign mem[556] = 12'd3539;
    assign mem[557] = 12'd3538;
    assign mem[558] = 12'd3537;
    assign mem[559] = 12'd3536;
    assign mem[560] = 12'd3535;
    assign mem[561] = 12'd3534;
    assign mem[562] = 12'd3533;
    assign mem[563] = 12'd3532;
    assign mem[564] = 12'd3531;
    assign mem[565] = 12'd3530;
    assign mem[566] = 12'd3529;
    assign mem[567] = 12'd3528;
    assign mem[568] = 12'd3527;
    assign mem[569] = 12'd3526;
    assign mem[570] = 12'd3525;
    assign mem[571] = 12'd3524;
    assign mem[572] = 12'd3523;
    assign mem[573] = 12'd3522;
    assign mem[574] = 12'd3521;
    assign mem[575] = 12'd3520;
    assign mem[576] = 12'd3519;
    assign mem[577] = 12'd3518;
    assign mem[578] = 12'd3517;
    assign mem[579] = 12'd3516;
    assign mem[580] = 12'd3515;
    assign mem[581] = 12'd3514;
    assign mem[582] = 12'd3513;
    assign mem[583] = 12'd3512;
    assign mem[584] = 12'd3511;
    assign mem[585] = 12'd3510;
    assign mem[586] = 12'd3509;
    assign mem[587] = 12'd3508;
    assign mem[588] = 12'd3507;
    assign mem[589] = 12'd3506;
    assign mem[590] = 12'd3505;
    assign mem[591] = 12'd3504;
    assign mem[592] = 12'd3503;
    assign mem[593] = 12'd3502;
    assign mem[594] = 12'd3501;
    assign mem[595] = 12'd3500;
    assign mem[596] = 12'd3499;
    assign mem[597] = 12'd3498;
    assign mem[598] = 12'd3497;
    assign mem[599] = 12'd3496;
    assign mem[600] = 12'd3495;
    assign mem[601] = 12'd3494;
    assign mem[602] = 12'd3493;
    assign mem[603] = 12'd3492;
    assign mem[604] = 12'd3491;
    assign mem[605] = 12'd3490;
    assign mem[606] = 12'd3489;
    assign mem[607] = 12'd3488;
    assign mem[608] = 12'd3487;
    assign mem[609] = 12'd3486;
    assign mem[610] = 12'd3485;
    assign mem[611] = 12'd3484;
    assign mem[612] = 12'd3483;
    assign mem[613] = 12'd3482;
    assign mem[614] = 12'd3481;
    assign mem[615] = 12'd3480;
    assign mem[616] = 12'd3479;
    assign mem[617] = 12'd3478;
    assign mem[618] = 12'd3477;
    assign mem[619] = 12'd3476;
    assign mem[620] = 12'd3475;
    assign mem[621] = 12'd3474;
    assign mem[622] = 12'd3473;
    assign mem[623] = 12'd3472;
    assign mem[624] = 12'd3471;
    assign mem[625] = 12'd3470;
    assign mem[626] = 12'd3469;
    assign mem[627] = 12'd3468;
    assign mem[628] = 12'd3467;
    assign mem[629] = 12'd3466;
    assign mem[630] = 12'd3465;
    assign mem[631] = 12'd3464;
    assign mem[632] = 12'd3463;
    assign mem[633] = 12'd3462;
    assign mem[634] = 12'd3461;
    assign mem[635] = 12'd3460;
    assign mem[636] = 12'd3459;
    assign mem[637] = 12'd3458;
    assign mem[638] = 12'd3457;
    assign mem[639] = 12'd3456;
    assign mem[640] = 12'd3455;
    assign mem[641] = 12'd3454;
    assign mem[642] = 12'd3453;
    assign mem[643] = 12'd3452;
    assign mem[644] = 12'd3451;
    assign mem[645] = 12'd3450;
    assign mem[646] = 12'd3449;
    assign mem[647] = 12'd3448;
    assign mem[648] = 12'd3447;
    assign mem[649] = 12'd3446;
    assign mem[650] = 12'd3445;
    assign mem[651] = 12'd3444;
    assign mem[652] = 12'd3443;
    assign mem[653] = 12'd3442;
    assign mem[654] = 12'd3441;
    assign mem[655] = 12'd3440;
    assign mem[656] = 12'd3439;
    assign mem[657] = 12'd3438;
    assign mem[658] = 12'd3437;
    assign mem[659] = 12'd3436;
    assign mem[660] = 12'd3435;
    assign mem[661] = 12'd3434;
    assign mem[662] = 12'd3433;
    assign mem[663] = 12'd3432;
    assign mem[664] = 12'd3431;
    assign mem[665] = 12'd3430;
    assign mem[666] = 12'd3429;
    assign mem[667] = 12'd3428;
    assign mem[668] = 12'd3427;
    assign mem[669] = 12'd3426;
    assign mem[670] = 12'd3425;
    assign mem[671] = 12'd3424;
    assign mem[672] = 12'd3423;
    assign mem[673] = 12'd3422;
    assign mem[674] = 12'd3421;
    assign mem[675] = 12'd3420;
    assign mem[676] = 12'd3419;
    assign mem[677] = 12'd3418;
    assign mem[678] = 12'd3417;
    assign mem[679] = 12'd3416;
    assign mem[680] = 12'd3415;
    assign mem[681] = 12'd3414;
    assign mem[682] = 12'd3413;
    assign mem[683] = 12'd3412;
    assign mem[684] = 12'd3411;
    assign mem[685] = 12'd3410;
    assign mem[686] = 12'd3409;
    assign mem[687] = 12'd3408;
    assign mem[688] = 12'd3407;
    assign mem[689] = 12'd3406;
    assign mem[690] = 12'd3405;
    assign mem[691] = 12'd3404;
    assign mem[692] = 12'd3403;
    assign mem[693] = 12'd3402;
    assign mem[694] = 12'd3401;
    assign mem[695] = 12'd3400;
    assign mem[696] = 12'd3399;
    assign mem[697] = 12'd3398;
    assign mem[698] = 12'd3397;
    assign mem[699] = 12'd3396;
    assign mem[700] = 12'd3395;
    assign mem[701] = 12'd3394;
    assign mem[702] = 12'd3393;
    assign mem[703] = 12'd3392;
    assign mem[704] = 12'd3391;
    assign mem[705] = 12'd3390;
    assign mem[706] = 12'd3389;
    assign mem[707] = 12'd3388;
    assign mem[708] = 12'd3387;
    assign mem[709] = 12'd3386;
    assign mem[710] = 12'd3385;
    assign mem[711] = 12'd3384;
    assign mem[712] = 12'd3383;
    assign mem[713] = 12'd3382;
    assign mem[714] = 12'd3381;
    assign mem[715] = 12'd3380;
    assign mem[716] = 12'd3379;
    assign mem[717] = 12'd3378;
    assign mem[718] = 12'd3377;
    assign mem[719] = 12'd3376;
    assign mem[720] = 12'd3375;
    assign mem[721] = 12'd3374;
    assign mem[722] = 12'd3373;
    assign mem[723] = 12'd3372;
    assign mem[724] = 12'd3371;
    assign mem[725] = 12'd3370;
    assign mem[726] = 12'd3369;
    assign mem[727] = 12'd3368;
    assign mem[728] = 12'd3367;
    assign mem[729] = 12'd3366;
    assign mem[730] = 12'd3365;
    assign mem[731] = 12'd3364;
    assign mem[732] = 12'd3363;
    assign mem[733] = 12'd3362;
    assign mem[734] = 12'd3361;
    assign mem[735] = 12'd3360;
    assign mem[736] = 12'd3359;
    assign mem[737] = 12'd3358;
    assign mem[738] = 12'd3357;
    assign mem[739] = 12'd3356;
    assign mem[740] = 12'd3355;
    assign mem[741] = 12'd3354;
    assign mem[742] = 12'd3353;
    assign mem[743] = 12'd3352;
    assign mem[744] = 12'd3351;
    assign mem[745] = 12'd3350;
    assign mem[746] = 12'd3349;
    assign mem[747] = 12'd3348;
    assign mem[748] = 12'd3347;
    assign mem[749] = 12'd3346;
    assign mem[750] = 12'd3345;
    assign mem[751] = 12'd3344;
    assign mem[752] = 12'd3343;
    assign mem[753] = 12'd3342;
    assign mem[754] = 12'd3341;
    assign mem[755] = 12'd3340;
    assign mem[756] = 12'd3339;
    assign mem[757] = 12'd3338;
    assign mem[758] = 12'd3337;
    assign mem[759] = 12'd3336;
    assign mem[760] = 12'd3335;
    assign mem[761] = 12'd3334;
    assign mem[762] = 12'd3333;
    assign mem[763] = 12'd3332;
    assign mem[764] = 12'd3331;
    assign mem[765] = 12'd3330;
    assign mem[766] = 12'd3329;
    assign mem[767] = 12'd3328;
    assign mem[768] = 12'd3327;
    assign mem[769] = 12'd3326;
    assign mem[770] = 12'd3325;
    assign mem[771] = 12'd3324;
    assign mem[772] = 12'd3323;
    assign mem[773] = 12'd3322;
    assign mem[774] = 12'd3321;
    assign mem[775] = 12'd3320;
    assign mem[776] = 12'd3319;
    assign mem[777] = 12'd3318;
    assign mem[778] = 12'd3317;
    assign mem[779] = 12'd3316;
    assign mem[780] = 12'd3315;
    assign mem[781] = 12'd3314;
    assign mem[782] = 12'd3313;
    assign mem[783] = 12'd3312;
    assign mem[784] = 12'd3311;
    assign mem[785] = 12'd3310;
    assign mem[786] = 12'd3309;
    assign mem[787] = 12'd3308;
    assign mem[788] = 12'd3307;
    assign mem[789] = 12'd3306;
    assign mem[790] = 12'd3305;
    assign mem[791] = 12'd3304;
    assign mem[792] = 12'd3303;
    assign mem[793] = 12'd3302;
    assign mem[794] = 12'd3301;
    assign mem[795] = 12'd3300;
    assign mem[796] = 12'd3299;
    assign mem[797] = 12'd3298;
    assign mem[798] = 12'd3297;
    assign mem[799] = 12'd3296;
    assign mem[800] = 12'd3295;
    assign mem[801] = 12'd3294;
    assign mem[802] = 12'd3293;
    assign mem[803] = 12'd3292;
    assign mem[804] = 12'd3291;
    assign mem[805] = 12'd3290;
    assign mem[806] = 12'd3289;
    assign mem[807] = 12'd3288;
    assign mem[808] = 12'd3287;
    assign mem[809] = 12'd3286;
    assign mem[810] = 12'd3285;
    assign mem[811] = 12'd3284;
    assign mem[812] = 12'd3283;
    assign mem[813] = 12'd3282;
    assign mem[814] = 12'd3281;
    assign mem[815] = 12'd3280;
    assign mem[816] = 12'd3279;
    assign mem[817] = 12'd3278;
    assign mem[818] = 12'd3277;
    assign mem[819] = 12'd3276;
    assign mem[820] = 12'd3275;
    assign mem[821] = 12'd3274;
    assign mem[822] = 12'd3273;
    assign mem[823] = 12'd3272;
    assign mem[824] = 12'd3271;
    assign mem[825] = 12'd3270;
    assign mem[826] = 12'd3269;
    assign mem[827] = 12'd3268;
    assign mem[828] = 12'd3267;
    assign mem[829] = 12'd3266;
    assign mem[830] = 12'd3265;
    assign mem[831] = 12'd3264;
    assign mem[832] = 12'd3263;
    assign mem[833] = 12'd3262;
    assign mem[834] = 12'd3261;
    assign mem[835] = 12'd3260;
    assign mem[836] = 12'd3259;
    assign mem[837] = 12'd3258;
    assign mem[838] = 12'd3257;
    assign mem[839] = 12'd3256;
    assign mem[840] = 12'd3255;
    assign mem[841] = 12'd3254;
    assign mem[842] = 12'd3253;
    assign mem[843] = 12'd3252;
    assign mem[844] = 12'd3251;
    assign mem[845] = 12'd3250;
    assign mem[846] = 12'd3249;
    assign mem[847] = 12'd3248;
    assign mem[848] = 12'd3247;
    assign mem[849] = 12'd3246;
    assign mem[850] = 12'd3245;
    assign mem[851] = 12'd3244;
    assign mem[852] = 12'd3243;
    assign mem[853] = 12'd3242;
    assign mem[854] = 12'd3241;
    assign mem[855] = 12'd3240;
    assign mem[856] = 12'd3239;
    assign mem[857] = 12'd3238;
    assign mem[858] = 12'd3237;
    assign mem[859] = 12'd3236;
    assign mem[860] = 12'd3235;
    assign mem[861] = 12'd3234;
    assign mem[862] = 12'd3233;
    assign mem[863] = 12'd3232;
    assign mem[864] = 12'd3231;
    assign mem[865] = 12'd3230;
    assign mem[866] = 12'd3229;
    assign mem[867] = 12'd3228;
    assign mem[868] = 12'd3227;
    assign mem[869] = 12'd3226;
    assign mem[870] = 12'd3225;
    assign mem[871] = 12'd3224;
    assign mem[872] = 12'd3223;
    assign mem[873] = 12'd3222;
    assign mem[874] = 12'd3221;
    assign mem[875] = 12'd3220;
    assign mem[876] = 12'd3219;
    assign mem[877] = 12'd3218;
    assign mem[878] = 12'd3217;
    assign mem[879] = 12'd3216;
    assign mem[880] = 12'd3215;
    assign mem[881] = 12'd3214;
    assign mem[882] = 12'd3213;
    assign mem[883] = 12'd3212;
    assign mem[884] = 12'd3211;
    assign mem[885] = 12'd3210;
    assign mem[886] = 12'd3209;
    assign mem[887] = 12'd3208;
    assign mem[888] = 12'd3207;
    assign mem[889] = 12'd3206;
    assign mem[890] = 12'd3205;
    assign mem[891] = 12'd3204;
    assign mem[892] = 12'd3203;
    assign mem[893] = 12'd3202;
    assign mem[894] = 12'd3201;
    assign mem[895] = 12'd3200;
    assign mem[896] = 12'd3199;
    assign mem[897] = 12'd3198;
    assign mem[898] = 12'd3197;
    assign mem[899] = 12'd3196;
    assign mem[900] = 12'd3195;
    assign mem[901] = 12'd3194;
    assign mem[902] = 12'd3193;
    assign mem[903] = 12'd3192;
    assign mem[904] = 12'd3191;
    assign mem[905] = 12'd3190;
    assign mem[906] = 12'd3189;
    assign mem[907] = 12'd3188;
    assign mem[908] = 12'd3187;
    assign mem[909] = 12'd3186;
    assign mem[910] = 12'd3185;
    assign mem[911] = 12'd3184;
    assign mem[912] = 12'd3183;
    assign mem[913] = 12'd3182;
    assign mem[914] = 12'd3181;
    assign mem[915] = 12'd3180;
    assign mem[916] = 12'd3179;
    assign mem[917] = 12'd3178;
    assign mem[918] = 12'd3177;
    assign mem[919] = 12'd3176;
    assign mem[920] = 12'd3175;
    assign mem[921] = 12'd3174;
    assign mem[922] = 12'd3173;
    assign mem[923] = 12'd3172;
    assign mem[924] = 12'd3171;
    assign mem[925] = 12'd3170;
    assign mem[926] = 12'd3169;
    assign mem[927] = 12'd3168;
    assign mem[928] = 12'd3167;
    assign mem[929] = 12'd3166;
    assign mem[930] = 12'd3165;
    assign mem[931] = 12'd3164;
    assign mem[932] = 12'd3163;
    assign mem[933] = 12'd3162;
    assign mem[934] = 12'd3161;
    assign mem[935] = 12'd3160;
    assign mem[936] = 12'd3159;
    assign mem[937] = 12'd3158;
    assign mem[938] = 12'd3157;
    assign mem[939] = 12'd3156;
    assign mem[940] = 12'd3155;
    assign mem[941] = 12'd3154;
    assign mem[942] = 12'd3153;
    assign mem[943] = 12'd3152;
    assign mem[944] = 12'd3151;
    assign mem[945] = 12'd3150;
    assign mem[946] = 12'd3149;
    assign mem[947] = 12'd3148;
    assign mem[948] = 12'd3147;
    assign mem[949] = 12'd3146;
    assign mem[950] = 12'd3145;
    assign mem[951] = 12'd3144;
    assign mem[952] = 12'd3143;
    assign mem[953] = 12'd3142;
    assign mem[954] = 12'd3141;
    assign mem[955] = 12'd3140;
    assign mem[956] = 12'd3139;
    assign mem[957] = 12'd3138;
    assign mem[958] = 12'd3137;
    assign mem[959] = 12'd3136;
    assign mem[960] = 12'd3135;
    assign mem[961] = 12'd3134;
    assign mem[962] = 12'd3133;
    assign mem[963] = 12'd3132;
    assign mem[964] = 12'd3131;
    assign mem[965] = 12'd3130;
    assign mem[966] = 12'd3129;
    assign mem[967] = 12'd3128;
    assign mem[968] = 12'd3127;
    assign mem[969] = 12'd3126;
    assign mem[970] = 12'd3125;
    assign mem[971] = 12'd3124;
    assign mem[972] = 12'd3123;
    assign mem[973] = 12'd3122;
    assign mem[974] = 12'd3121;
    assign mem[975] = 12'd3120;
    assign mem[976] = 12'd3119;
    assign mem[977] = 12'd3118;
    assign mem[978] = 12'd3117;
    assign mem[979] = 12'd3116;
    assign mem[980] = 12'd3115;
    assign mem[981] = 12'd3114;
    assign mem[982] = 12'd3113;
    assign mem[983] = 12'd3112;
    assign mem[984] = 12'd3111;
    assign mem[985] = 12'd3110;
    assign mem[986] = 12'd3109;
    assign mem[987] = 12'd3108;
    assign mem[988] = 12'd3107;
    assign mem[989] = 12'd3106;
    assign mem[990] = 12'd3105;
    assign mem[991] = 12'd3104;
    assign mem[992] = 12'd3103;
    assign mem[993] = 12'd3102;
    assign mem[994] = 12'd3101;
    assign mem[995] = 12'd3100;
    assign mem[996] = 12'd3099;
    assign mem[997] = 12'd3098;
    assign mem[998] = 12'd3097;
    assign mem[999] = 12'd3096;
    assign mem[1000] = 12'd3095;
    assign mem[1001] = 12'd3094;
    assign mem[1002] = 12'd3093;
    assign mem[1003] = 12'd3092;
    assign mem[1004] = 12'd3091;
    assign mem[1005] = 12'd3090;
    assign mem[1006] = 12'd3089;
    assign mem[1007] = 12'd3088;
    assign mem[1008] = 12'd3087;
    assign mem[1009] = 12'd3086;
    assign mem[1010] = 12'd3085;
    assign mem[1011] = 12'd3084;
    assign mem[1012] = 12'd3083;
    assign mem[1013] = 12'd3082;
    assign mem[1014] = 12'd3081;
    assign mem[1015] = 12'd3080;
    assign mem[1016] = 12'd3079;
    assign mem[1017] = 12'd3078;
    assign mem[1018] = 12'd3077;
    assign mem[1019] = 12'd3076;
    assign mem[1020] = 12'd3075;
    assign mem[1021] = 12'd3074;
    assign mem[1022] = 12'd3073;
    assign mem[1023] = 12'd3072;
    assign mem[1024] = 12'd3071;
    assign mem[1025] = 12'd3070;
    assign mem[1026] = 12'd3069;
    assign mem[1027] = 12'd3068;
    assign mem[1028] = 12'd3067;
    assign mem[1029] = 12'd3066;
    assign mem[1030] = 12'd3065;
    assign mem[1031] = 12'd3064;
    assign mem[1032] = 12'd3063;
    assign mem[1033] = 12'd3062;
    assign mem[1034] = 12'd3061;
    assign mem[1035] = 12'd3060;
    assign mem[1036] = 12'd3059;
    assign mem[1037] = 12'd3058;
    assign mem[1038] = 12'd3057;
    assign mem[1039] = 12'd3056;
    assign mem[1040] = 12'd3055;
    assign mem[1041] = 12'd3054;
    assign mem[1042] = 12'd3053;
    assign mem[1043] = 12'd3052;
    assign mem[1044] = 12'd3051;
    assign mem[1045] = 12'd3050;
    assign mem[1046] = 12'd3049;
    assign mem[1047] = 12'd3048;
    assign mem[1048] = 12'd3047;
    assign mem[1049] = 12'd3046;
    assign mem[1050] = 12'd3045;
    assign mem[1051] = 12'd3044;
    assign mem[1052] = 12'd3043;
    assign mem[1053] = 12'd3042;
    assign mem[1054] = 12'd3041;
    assign mem[1055] = 12'd3040;
    assign mem[1056] = 12'd3039;
    assign mem[1057] = 12'd3038;
    assign mem[1058] = 12'd3037;
    assign mem[1059] = 12'd3036;
    assign mem[1060] = 12'd3035;
    assign mem[1061] = 12'd3034;
    assign mem[1062] = 12'd3033;
    assign mem[1063] = 12'd3032;
    assign mem[1064] = 12'd3031;
    assign mem[1065] = 12'd3030;
    assign mem[1066] = 12'd3029;
    assign mem[1067] = 12'd3028;
    assign mem[1068] = 12'd3027;
    assign mem[1069] = 12'd3026;
    assign mem[1070] = 12'd3025;
    assign mem[1071] = 12'd3024;
    assign mem[1072] = 12'd3023;
    assign mem[1073] = 12'd3022;
    assign mem[1074] = 12'd3021;
    assign mem[1075] = 12'd3020;
    assign mem[1076] = 12'd3019;
    assign mem[1077] = 12'd3018;
    assign mem[1078] = 12'd3017;
    assign mem[1079] = 12'd3016;
    assign mem[1080] = 12'd3015;
    assign mem[1081] = 12'd3014;
    assign mem[1082] = 12'd3013;
    assign mem[1083] = 12'd3012;
    assign mem[1084] = 12'd3011;
    assign mem[1085] = 12'd3010;
    assign mem[1086] = 12'd3009;
    assign mem[1087] = 12'd3008;
    assign mem[1088] = 12'd3007;
    assign mem[1089] = 12'd3006;
    assign mem[1090] = 12'd3005;
    assign mem[1091] = 12'd3004;
    assign mem[1092] = 12'd3003;
    assign mem[1093] = 12'd3002;
    assign mem[1094] = 12'd3001;
    assign mem[1095] = 12'd3000;
    assign mem[1096] = 12'd2999;
    assign mem[1097] = 12'd2998;
    assign mem[1098] = 12'd2997;
    assign mem[1099] = 12'd2996;
    assign mem[1100] = 12'd2995;
    assign mem[1101] = 12'd2994;
    assign mem[1102] = 12'd2993;
    assign mem[1103] = 12'd2992;
    assign mem[1104] = 12'd2991;
    assign mem[1105] = 12'd2990;
    assign mem[1106] = 12'd2989;
    assign mem[1107] = 12'd2988;
    assign mem[1108] = 12'd2987;
    assign mem[1109] = 12'd2986;
    assign mem[1110] = 12'd2985;
    assign mem[1111] = 12'd2984;
    assign mem[1112] = 12'd2983;
    assign mem[1113] = 12'd2982;
    assign mem[1114] = 12'd2981;
    assign mem[1115] = 12'd2980;
    assign mem[1116] = 12'd2979;
    assign mem[1117] = 12'd2978;
    assign mem[1118] = 12'd2977;
    assign mem[1119] = 12'd2976;
    assign mem[1120] = 12'd2975;
    assign mem[1121] = 12'd2974;
    assign mem[1122] = 12'd2973;
    assign mem[1123] = 12'd2972;
    assign mem[1124] = 12'd2971;
    assign mem[1125] = 12'd2970;
    assign mem[1126] = 12'd2969;
    assign mem[1127] = 12'd2968;
    assign mem[1128] = 12'd2967;
    assign mem[1129] = 12'd2966;
    assign mem[1130] = 12'd2965;
    assign mem[1131] = 12'd2964;
    assign mem[1132] = 12'd2963;
    assign mem[1133] = 12'd2962;
    assign mem[1134] = 12'd2961;
    assign mem[1135] = 12'd2960;
    assign mem[1136] = 12'd2959;
    assign mem[1137] = 12'd2958;
    assign mem[1138] = 12'd2957;
    assign mem[1139] = 12'd2956;
    assign mem[1140] = 12'd2955;
    assign mem[1141] = 12'd2954;
    assign mem[1142] = 12'd2953;
    assign mem[1143] = 12'd2952;
    assign mem[1144] = 12'd2951;
    assign mem[1145] = 12'd2950;
    assign mem[1146] = 12'd2949;
    assign mem[1147] = 12'd2948;
    assign mem[1148] = 12'd2947;
    assign mem[1149] = 12'd2946;
    assign mem[1150] = 12'd2945;
    assign mem[1151] = 12'd2944;
    assign mem[1152] = 12'd2943;
    assign mem[1153] = 12'd2942;
    assign mem[1154] = 12'd2941;
    assign mem[1155] = 12'd2940;
    assign mem[1156] = 12'd2939;
    assign mem[1157] = 12'd2938;
    assign mem[1158] = 12'd2937;
    assign mem[1159] = 12'd2936;
    assign mem[1160] = 12'd2935;
    assign mem[1161] = 12'd2934;
    assign mem[1162] = 12'd2933;
    assign mem[1163] = 12'd2932;
    assign mem[1164] = 12'd2931;
    assign mem[1165] = 12'd2930;
    assign mem[1166] = 12'd2929;
    assign mem[1167] = 12'd2928;
    assign mem[1168] = 12'd2927;
    assign mem[1169] = 12'd2926;
    assign mem[1170] = 12'd2925;
    assign mem[1171] = 12'd2924;
    assign mem[1172] = 12'd2923;
    assign mem[1173] = 12'd2922;
    assign mem[1174] = 12'd2921;
    assign mem[1175] = 12'd2920;
    assign mem[1176] = 12'd2919;
    assign mem[1177] = 12'd2918;
    assign mem[1178] = 12'd2917;
    assign mem[1179] = 12'd2916;
    assign mem[1180] = 12'd2915;
    assign mem[1181] = 12'd2914;
    assign mem[1182] = 12'd2913;
    assign mem[1183] = 12'd2912;
    assign mem[1184] = 12'd2911;
    assign mem[1185] = 12'd2910;
    assign mem[1186] = 12'd2909;
    assign mem[1187] = 12'd2908;
    assign mem[1188] = 12'd2907;
    assign mem[1189] = 12'd2906;
    assign mem[1190] = 12'd2905;
    assign mem[1191] = 12'd2904;
    assign mem[1192] = 12'd2903;
    assign mem[1193] = 12'd2902;
    assign mem[1194] = 12'd2901;
    assign mem[1195] = 12'd2900;
    assign mem[1196] = 12'd2899;
    assign mem[1197] = 12'd2898;
    assign mem[1198] = 12'd2897;
    assign mem[1199] = 12'd2896;
    assign mem[1200] = 12'd2895;
    assign mem[1201] = 12'd2894;
    assign mem[1202] = 12'd2893;
    assign mem[1203] = 12'd2892;
    assign mem[1204] = 12'd2891;
    assign mem[1205] = 12'd2890;
    assign mem[1206] = 12'd2889;
    assign mem[1207] = 12'd2888;
    assign mem[1208] = 12'd2887;
    assign mem[1209] = 12'd2886;
    assign mem[1210] = 12'd2885;
    assign mem[1211] = 12'd2884;
    assign mem[1212] = 12'd2883;
    assign mem[1213] = 12'd2882;
    assign mem[1214] = 12'd2881;
    assign mem[1215] = 12'd2880;
    assign mem[1216] = 12'd2879;
    assign mem[1217] = 12'd2878;
    assign mem[1218] = 12'd2877;
    assign mem[1219] = 12'd2876;
    assign mem[1220] = 12'd2875;
    assign mem[1221] = 12'd2874;
    assign mem[1222] = 12'd2873;
    assign mem[1223] = 12'd2872;
    assign mem[1224] = 12'd2871;
    assign mem[1225] = 12'd2870;
    assign mem[1226] = 12'd2869;
    assign mem[1227] = 12'd2868;
    assign mem[1228] = 12'd2867;
    assign mem[1229] = 12'd2866;
    assign mem[1230] = 12'd2865;
    assign mem[1231] = 12'd2864;
    assign mem[1232] = 12'd2863;
    assign mem[1233] = 12'd2862;
    assign mem[1234] = 12'd2861;
    assign mem[1235] = 12'd2860;
    assign mem[1236] = 12'd2859;
    assign mem[1237] = 12'd2858;
    assign mem[1238] = 12'd2857;
    assign mem[1239] = 12'd2856;
    assign mem[1240] = 12'd2855;
    assign mem[1241] = 12'd2854;
    assign mem[1242] = 12'd2853;
    assign mem[1243] = 12'd2852;
    assign mem[1244] = 12'd2851;
    assign mem[1245] = 12'd2850;
    assign mem[1246] = 12'd2849;
    assign mem[1247] = 12'd2848;
    assign mem[1248] = 12'd2847;
    assign mem[1249] = 12'd2846;
    assign mem[1250] = 12'd2845;
    assign mem[1251] = 12'd2844;
    assign mem[1252] = 12'd2843;
    assign mem[1253] = 12'd2842;
    assign mem[1254] = 12'd2841;
    assign mem[1255] = 12'd2840;
    assign mem[1256] = 12'd2839;
    assign mem[1257] = 12'd2838;
    assign mem[1258] = 12'd2837;
    assign mem[1259] = 12'd2836;
    assign mem[1260] = 12'd2835;
    assign mem[1261] = 12'd2834;
    assign mem[1262] = 12'd2833;
    assign mem[1263] = 12'd2832;
    assign mem[1264] = 12'd2831;
    assign mem[1265] = 12'd2830;
    assign mem[1266] = 12'd2829;
    assign mem[1267] = 12'd2828;
    assign mem[1268] = 12'd2827;
    assign mem[1269] = 12'd2826;
    assign mem[1270] = 12'd2825;
    assign mem[1271] = 12'd2824;
    assign mem[1272] = 12'd2823;
    assign mem[1273] = 12'd2822;
    assign mem[1274] = 12'd2821;
    assign mem[1275] = 12'd2820;
    assign mem[1276] = 12'd2819;
    assign mem[1277] = 12'd2818;
    assign mem[1278] = 12'd2817;
    assign mem[1279] = 12'd2816;
    assign mem[1280] = 12'd2815;
    assign mem[1281] = 12'd2814;
    assign mem[1282] = 12'd2813;
    assign mem[1283] = 12'd2812;
    assign mem[1284] = 12'd2811;
    assign mem[1285] = 12'd2810;
    assign mem[1286] = 12'd2809;
    assign mem[1287] = 12'd2808;
    assign mem[1288] = 12'd2807;
    assign mem[1289] = 12'd2806;
    assign mem[1290] = 12'd2805;
    assign mem[1291] = 12'd2804;
    assign mem[1292] = 12'd2803;
    assign mem[1293] = 12'd2802;
    assign mem[1294] = 12'd2801;
    assign mem[1295] = 12'd2800;
    assign mem[1296] = 12'd2799;
    assign mem[1297] = 12'd2798;
    assign mem[1298] = 12'd2797;
    assign mem[1299] = 12'd2796;
    assign mem[1300] = 12'd2795;
    assign mem[1301] = 12'd2794;
    assign mem[1302] = 12'd2793;
    assign mem[1303] = 12'd2792;
    assign mem[1304] = 12'd2791;
    assign mem[1305] = 12'd2790;
    assign mem[1306] = 12'd2789;
    assign mem[1307] = 12'd2788;
    assign mem[1308] = 12'd2787;
    assign mem[1309] = 12'd2786;
    assign mem[1310] = 12'd2785;
    assign mem[1311] = 12'd2784;
    assign mem[1312] = 12'd2783;
    assign mem[1313] = 12'd2782;
    assign mem[1314] = 12'd2781;
    assign mem[1315] = 12'd2780;
    assign mem[1316] = 12'd2779;
    assign mem[1317] = 12'd2778;
    assign mem[1318] = 12'd2777;
    assign mem[1319] = 12'd2776;
    assign mem[1320] = 12'd2775;
    assign mem[1321] = 12'd2774;
    assign mem[1322] = 12'd2773;
    assign mem[1323] = 12'd2772;
    assign mem[1324] = 12'd2771;
    assign mem[1325] = 12'd2770;
    assign mem[1326] = 12'd2769;
    assign mem[1327] = 12'd2768;
    assign mem[1328] = 12'd2767;
    assign mem[1329] = 12'd2766;
    assign mem[1330] = 12'd2765;
    assign mem[1331] = 12'd2764;
    assign mem[1332] = 12'd2763;
    assign mem[1333] = 12'd2762;
    assign mem[1334] = 12'd2761;
    assign mem[1335] = 12'd2760;
    assign mem[1336] = 12'd2759;
    assign mem[1337] = 12'd2758;
    assign mem[1338] = 12'd2757;
    assign mem[1339] = 12'd2756;
    assign mem[1340] = 12'd2755;
    assign mem[1341] = 12'd2754;
    assign mem[1342] = 12'd2753;
    assign mem[1343] = 12'd2752;
    assign mem[1344] = 12'd2751;
    assign mem[1345] = 12'd2750;
    assign mem[1346] = 12'd2749;
    assign mem[1347] = 12'd2748;
    assign mem[1348] = 12'd2747;
    assign mem[1349] = 12'd2746;
    assign mem[1350] = 12'd2745;
    assign mem[1351] = 12'd2744;
    assign mem[1352] = 12'd2743;
    assign mem[1353] = 12'd2742;
    assign mem[1354] = 12'd2741;
    assign mem[1355] = 12'd2740;
    assign mem[1356] = 12'd2739;
    assign mem[1357] = 12'd2738;
    assign mem[1358] = 12'd2737;
    assign mem[1359] = 12'd2736;
    assign mem[1360] = 12'd2735;
    assign mem[1361] = 12'd2734;
    assign mem[1362] = 12'd2733;
    assign mem[1363] = 12'd2732;
    assign mem[1364] = 12'd2731;
    assign mem[1365] = 12'd2730;
    assign mem[1366] = 12'd2729;
    assign mem[1367] = 12'd2728;
    assign mem[1368] = 12'd2727;
    assign mem[1369] = 12'd2726;
    assign mem[1370] = 12'd2725;
    assign mem[1371] = 12'd2724;
    assign mem[1372] = 12'd2723;
    assign mem[1373] = 12'd2722;
    assign mem[1374] = 12'd2721;
    assign mem[1375] = 12'd2720;
    assign mem[1376] = 12'd2719;
    assign mem[1377] = 12'd2718;
    assign mem[1378] = 12'd2717;
    assign mem[1379] = 12'd2716;
    assign mem[1380] = 12'd2715;
    assign mem[1381] = 12'd2714;
    assign mem[1382] = 12'd2713;
    assign mem[1383] = 12'd2712;
    assign mem[1384] = 12'd2711;
    assign mem[1385] = 12'd2710;
    assign mem[1386] = 12'd2709;
    assign mem[1387] = 12'd2708;
    assign mem[1388] = 12'd2707;
    assign mem[1389] = 12'd2706;
    assign mem[1390] = 12'd2705;
    assign mem[1391] = 12'd2704;
    assign mem[1392] = 12'd2703;
    assign mem[1393] = 12'd2702;
    assign mem[1394] = 12'd2701;
    assign mem[1395] = 12'd2700;
    assign mem[1396] = 12'd2699;
    assign mem[1397] = 12'd2698;
    assign mem[1398] = 12'd2697;
    assign mem[1399] = 12'd2696;
    assign mem[1400] = 12'd2695;
    assign mem[1401] = 12'd2694;
    assign mem[1402] = 12'd2693;
    assign mem[1403] = 12'd2692;
    assign mem[1404] = 12'd2691;
    assign mem[1405] = 12'd2690;
    assign mem[1406] = 12'd2689;
    assign mem[1407] = 12'd2688;
    assign mem[1408] = 12'd2687;
    assign mem[1409] = 12'd2686;
    assign mem[1410] = 12'd2685;
    assign mem[1411] = 12'd2684;
    assign mem[1412] = 12'd2683;
    assign mem[1413] = 12'd2682;
    assign mem[1414] = 12'd2681;
    assign mem[1415] = 12'd2680;
    assign mem[1416] = 12'd2679;
    assign mem[1417] = 12'd2678;
    assign mem[1418] = 12'd2677;
    assign mem[1419] = 12'd2676;
    assign mem[1420] = 12'd2675;
    assign mem[1421] = 12'd2674;
    assign mem[1422] = 12'd2673;
    assign mem[1423] = 12'd2672;
    assign mem[1424] = 12'd2671;
    assign mem[1425] = 12'd2670;
    assign mem[1426] = 12'd2669;
    assign mem[1427] = 12'd2668;
    assign mem[1428] = 12'd2667;
    assign mem[1429] = 12'd2666;
    assign mem[1430] = 12'd2665;
    assign mem[1431] = 12'd2664;
    assign mem[1432] = 12'd2663;
    assign mem[1433] = 12'd2662;
    assign mem[1434] = 12'd2661;
    assign mem[1435] = 12'd2660;
    assign mem[1436] = 12'd2659;
    assign mem[1437] = 12'd2658;
    assign mem[1438] = 12'd2657;
    assign mem[1439] = 12'd2656;
    assign mem[1440] = 12'd2655;
    assign mem[1441] = 12'd2654;
    assign mem[1442] = 12'd2653;
    assign mem[1443] = 12'd2652;
    assign mem[1444] = 12'd2651;
    assign mem[1445] = 12'd2650;
    assign mem[1446] = 12'd2649;
    assign mem[1447] = 12'd2648;
    assign mem[1448] = 12'd2647;
    assign mem[1449] = 12'd2646;
    assign mem[1450] = 12'd2645;
    assign mem[1451] = 12'd2644;
    assign mem[1452] = 12'd2643;
    assign mem[1453] = 12'd2642;
    assign mem[1454] = 12'd2641;
    assign mem[1455] = 12'd2640;
    assign mem[1456] = 12'd2639;
    assign mem[1457] = 12'd2638;
    assign mem[1458] = 12'd2637;
    assign mem[1459] = 12'd2636;
    assign mem[1460] = 12'd2635;
    assign mem[1461] = 12'd2634;
    assign mem[1462] = 12'd2633;
    assign mem[1463] = 12'd2632;
    assign mem[1464] = 12'd2631;
    assign mem[1465] = 12'd2630;
    assign mem[1466] = 12'd2629;
    assign mem[1467] = 12'd2628;
    assign mem[1468] = 12'd2627;
    assign mem[1469] = 12'd2626;
    assign mem[1470] = 12'd2625;
    assign mem[1471] = 12'd2624;
    assign mem[1472] = 12'd2623;
    assign mem[1473] = 12'd2622;
    assign mem[1474] = 12'd2621;
    assign mem[1475] = 12'd2620;
    assign mem[1476] = 12'd2619;
    assign mem[1477] = 12'd2618;
    assign mem[1478] = 12'd2617;
    assign mem[1479] = 12'd2616;
    assign mem[1480] = 12'd2615;
    assign mem[1481] = 12'd2614;
    assign mem[1482] = 12'd2613;
    assign mem[1483] = 12'd2612;
    assign mem[1484] = 12'd2611;
    assign mem[1485] = 12'd2610;
    assign mem[1486] = 12'd2609;
    assign mem[1487] = 12'd2608;
    assign mem[1488] = 12'd2607;
    assign mem[1489] = 12'd2606;
    assign mem[1490] = 12'd2605;
    assign mem[1491] = 12'd2604;
    assign mem[1492] = 12'd2603;
    assign mem[1493] = 12'd2602;
    assign mem[1494] = 12'd2601;
    assign mem[1495] = 12'd2600;
    assign mem[1496] = 12'd2599;
    assign mem[1497] = 12'd2598;
    assign mem[1498] = 12'd2597;
    assign mem[1499] = 12'd2596;
    assign mem[1500] = 12'd2595;
    assign mem[1501] = 12'd2594;
    assign mem[1502] = 12'd2593;
    assign mem[1503] = 12'd2592;
    assign mem[1504] = 12'd2591;
    assign mem[1505] = 12'd2590;
    assign mem[1506] = 12'd2589;
    assign mem[1507] = 12'd2588;
    assign mem[1508] = 12'd2587;
    assign mem[1509] = 12'd2586;
    assign mem[1510] = 12'd2585;
    assign mem[1511] = 12'd2584;
    assign mem[1512] = 12'd2583;
    assign mem[1513] = 12'd2582;
    assign mem[1514] = 12'd2581;
    assign mem[1515] = 12'd2580;
    assign mem[1516] = 12'd2579;
    assign mem[1517] = 12'd2578;
    assign mem[1518] = 12'd2577;
    assign mem[1519] = 12'd2576;
    assign mem[1520] = 12'd2575;
    assign mem[1521] = 12'd2574;
    assign mem[1522] = 12'd2573;
    assign mem[1523] = 12'd2572;
    assign mem[1524] = 12'd2571;
    assign mem[1525] = 12'd2570;
    assign mem[1526] = 12'd2569;
    assign mem[1527] = 12'd2568;
    assign mem[1528] = 12'd2567;
    assign mem[1529] = 12'd2566;
    assign mem[1530] = 12'd2565;
    assign mem[1531] = 12'd2564;
    assign mem[1532] = 12'd2563;
    assign mem[1533] = 12'd2562;
    assign mem[1534] = 12'd2561;
    assign mem[1535] = 12'd2560;
    assign mem[1536] = 12'd2559;
    assign mem[1537] = 12'd2558;
    assign mem[1538] = 12'd2557;
    assign mem[1539] = 12'd2556;
    assign mem[1540] = 12'd2555;
    assign mem[1541] = 12'd2554;
    assign mem[1542] = 12'd2553;
    assign mem[1543] = 12'd2552;
    assign mem[1544] = 12'd2551;
    assign mem[1545] = 12'd2550;
    assign mem[1546] = 12'd2549;
    assign mem[1547] = 12'd2548;
    assign mem[1548] = 12'd2547;
    assign mem[1549] = 12'd2546;
    assign mem[1550] = 12'd2545;
    assign mem[1551] = 12'd2544;
    assign mem[1552] = 12'd2543;
    assign mem[1553] = 12'd2542;
    assign mem[1554] = 12'd2541;
    assign mem[1555] = 12'd2540;
    assign mem[1556] = 12'd2539;
    assign mem[1557] = 12'd2538;
    assign mem[1558] = 12'd2537;
    assign mem[1559] = 12'd2536;
    assign mem[1560] = 12'd2535;
    assign mem[1561] = 12'd2534;
    assign mem[1562] = 12'd2533;
    assign mem[1563] = 12'd2532;
    assign mem[1564] = 12'd2531;
    assign mem[1565] = 12'd2530;
    assign mem[1566] = 12'd2529;
    assign mem[1567] = 12'd2528;
    assign mem[1568] = 12'd2527;
    assign mem[1569] = 12'd2526;
    assign mem[1570] = 12'd2525;
    assign mem[1571] = 12'd2524;
    assign mem[1572] = 12'd2523;
    assign mem[1573] = 12'd2522;
    assign mem[1574] = 12'd2521;
    assign mem[1575] = 12'd2520;
    assign mem[1576] = 12'd2519;
    assign mem[1577] = 12'd2518;
    assign mem[1578] = 12'd2517;
    assign mem[1579] = 12'd2516;
    assign mem[1580] = 12'd2515;
    assign mem[1581] = 12'd2514;
    assign mem[1582] = 12'd2513;
    assign mem[1583] = 12'd2512;
    assign mem[1584] = 12'd2511;
    assign mem[1585] = 12'd2510;
    assign mem[1586] = 12'd2509;
    assign mem[1587] = 12'd2508;
    assign mem[1588] = 12'd2507;
    assign mem[1589] = 12'd2506;
    assign mem[1590] = 12'd2505;
    assign mem[1591] = 12'd2504;
    assign mem[1592] = 12'd2503;
    assign mem[1593] = 12'd2502;
    assign mem[1594] = 12'd2501;
    assign mem[1595] = 12'd2500;
    assign mem[1596] = 12'd2499;
    assign mem[1597] = 12'd2498;
    assign mem[1598] = 12'd2497;
    assign mem[1599] = 12'd2496;
    assign mem[1600] = 12'd2495;
    assign mem[1601] = 12'd2494;
    assign mem[1602] = 12'd2493;
    assign mem[1603] = 12'd2492;
    assign mem[1604] = 12'd2491;
    assign mem[1605] = 12'd2490;
    assign mem[1606] = 12'd2489;
    assign mem[1607] = 12'd2488;
    assign mem[1608] = 12'd2487;
    assign mem[1609] = 12'd2486;
    assign mem[1610] = 12'd2485;
    assign mem[1611] = 12'd2484;
    assign mem[1612] = 12'd2483;
    assign mem[1613] = 12'd2482;
    assign mem[1614] = 12'd2481;
    assign mem[1615] = 12'd2480;
    assign mem[1616] = 12'd2479;
    assign mem[1617] = 12'd2478;
    assign mem[1618] = 12'd2477;
    assign mem[1619] = 12'd2476;
    assign mem[1620] = 12'd2475;
    assign mem[1621] = 12'd2474;
    assign mem[1622] = 12'd2473;
    assign mem[1623] = 12'd2472;
    assign mem[1624] = 12'd2471;
    assign mem[1625] = 12'd2470;
    assign mem[1626] = 12'd2469;
    assign mem[1627] = 12'd2468;
    assign mem[1628] = 12'd2467;
    assign mem[1629] = 12'd2466;
    assign mem[1630] = 12'd2465;
    assign mem[1631] = 12'd2464;
    assign mem[1632] = 12'd2463;
    assign mem[1633] = 12'd2462;
    assign mem[1634] = 12'd2461;
    assign mem[1635] = 12'd2460;
    assign mem[1636] = 12'd2459;
    assign mem[1637] = 12'd2458;
    assign mem[1638] = 12'd2457;
    assign mem[1639] = 12'd2456;
    assign mem[1640] = 12'd2455;
    assign mem[1641] = 12'd2454;
    assign mem[1642] = 12'd2453;
    assign mem[1643] = 12'd2452;
    assign mem[1644] = 12'd2451;
    assign mem[1645] = 12'd2450;
    assign mem[1646] = 12'd2449;
    assign mem[1647] = 12'd2448;
    assign mem[1648] = 12'd2447;
    assign mem[1649] = 12'd2446;
    assign mem[1650] = 12'd2445;
    assign mem[1651] = 12'd2444;
    assign mem[1652] = 12'd2443;
    assign mem[1653] = 12'd2442;
    assign mem[1654] = 12'd2441;
    assign mem[1655] = 12'd2440;
    assign mem[1656] = 12'd2439;
    assign mem[1657] = 12'd2438;
    assign mem[1658] = 12'd2437;
    assign mem[1659] = 12'd2436;
    assign mem[1660] = 12'd2435;
    assign mem[1661] = 12'd2434;
    assign mem[1662] = 12'd2433;
    assign mem[1663] = 12'd2432;
    assign mem[1664] = 12'd2431;
    assign mem[1665] = 12'd2430;
    assign mem[1666] = 12'd2429;
    assign mem[1667] = 12'd2428;
    assign mem[1668] = 12'd2427;
    assign mem[1669] = 12'd2426;
    assign mem[1670] = 12'd2425;
    assign mem[1671] = 12'd2424;
    assign mem[1672] = 12'd2423;
    assign mem[1673] = 12'd2422;
    assign mem[1674] = 12'd2421;
    assign mem[1675] = 12'd2420;
    assign mem[1676] = 12'd2419;
    assign mem[1677] = 12'd2418;
    assign mem[1678] = 12'd2417;
    assign mem[1679] = 12'd2416;
    assign mem[1680] = 12'd2415;
    assign mem[1681] = 12'd2414;
    assign mem[1682] = 12'd2413;
    assign mem[1683] = 12'd2412;
    assign mem[1684] = 12'd2411;
    assign mem[1685] = 12'd2410;
    assign mem[1686] = 12'd2409;
    assign mem[1687] = 12'd2408;
    assign mem[1688] = 12'd2407;
    assign mem[1689] = 12'd2406;
    assign mem[1690] = 12'd2405;
    assign mem[1691] = 12'd2404;
    assign mem[1692] = 12'd2403;
    assign mem[1693] = 12'd2402;
    assign mem[1694] = 12'd2401;
    assign mem[1695] = 12'd2400;
    assign mem[1696] = 12'd2399;
    assign mem[1697] = 12'd2398;
    assign mem[1698] = 12'd2397;
    assign mem[1699] = 12'd2396;
    assign mem[1700] = 12'd2395;
    assign mem[1701] = 12'd2394;
    assign mem[1702] = 12'd2393;
    assign mem[1703] = 12'd2392;
    assign mem[1704] = 12'd2391;
    assign mem[1705] = 12'd2390;
    assign mem[1706] = 12'd2389;
    assign mem[1707] = 12'd2388;
    assign mem[1708] = 12'd2387;
    assign mem[1709] = 12'd2386;
    assign mem[1710] = 12'd2385;
    assign mem[1711] = 12'd2384;
    assign mem[1712] = 12'd2383;
    assign mem[1713] = 12'd2382;
    assign mem[1714] = 12'd2381;
    assign mem[1715] = 12'd2380;
    assign mem[1716] = 12'd2379;
    assign mem[1717] = 12'd2378;
    assign mem[1718] = 12'd2377;
    assign mem[1719] = 12'd2376;
    assign mem[1720] = 12'd2375;
    assign mem[1721] = 12'd2374;
    assign mem[1722] = 12'd2373;
    assign mem[1723] = 12'd2372;
    assign mem[1724] = 12'd2371;
    assign mem[1725] = 12'd2370;
    assign mem[1726] = 12'd2369;
    assign mem[1727] = 12'd2368;
    assign mem[1728] = 12'd2367;
    assign mem[1729] = 12'd2366;
    assign mem[1730] = 12'd2365;
    assign mem[1731] = 12'd2364;
    assign mem[1732] = 12'd2363;
    assign mem[1733] = 12'd2362;
    assign mem[1734] = 12'd2361;
    assign mem[1735] = 12'd2360;
    assign mem[1736] = 12'd2359;
    assign mem[1737] = 12'd2358;
    assign mem[1738] = 12'd2357;
    assign mem[1739] = 12'd2356;
    assign mem[1740] = 12'd2355;
    assign mem[1741] = 12'd2354;
    assign mem[1742] = 12'd2353;
    assign mem[1743] = 12'd2352;
    assign mem[1744] = 12'd2351;
    assign mem[1745] = 12'd2350;
    assign mem[1746] = 12'd2349;
    assign mem[1747] = 12'd2348;
    assign mem[1748] = 12'd2347;
    assign mem[1749] = 12'd2346;
    assign mem[1750] = 12'd2345;
    assign mem[1751] = 12'd2344;
    assign mem[1752] = 12'd2343;
    assign mem[1753] = 12'd2342;
    assign mem[1754] = 12'd2341;
    assign mem[1755] = 12'd2340;
    assign mem[1756] = 12'd2339;
    assign mem[1757] = 12'd2338;
    assign mem[1758] = 12'd2337;
    assign mem[1759] = 12'd2336;
    assign mem[1760] = 12'd2335;
    assign mem[1761] = 12'd2334;
    assign mem[1762] = 12'd2333;
    assign mem[1763] = 12'd2332;
    assign mem[1764] = 12'd2331;
    assign mem[1765] = 12'd2330;
    assign mem[1766] = 12'd2329;
    assign mem[1767] = 12'd2328;
    assign mem[1768] = 12'd2327;
    assign mem[1769] = 12'd2326;
    assign mem[1770] = 12'd2325;
    assign mem[1771] = 12'd2324;
    assign mem[1772] = 12'd2323;
    assign mem[1773] = 12'd2322;
    assign mem[1774] = 12'd2321;
    assign mem[1775] = 12'd2320;
    assign mem[1776] = 12'd2319;
    assign mem[1777] = 12'd2318;
    assign mem[1778] = 12'd2317;
    assign mem[1779] = 12'd2316;
    assign mem[1780] = 12'd2315;
    assign mem[1781] = 12'd2314;
    assign mem[1782] = 12'd2313;
    assign mem[1783] = 12'd2312;
    assign mem[1784] = 12'd2311;
    assign mem[1785] = 12'd2310;
    assign mem[1786] = 12'd2309;
    assign mem[1787] = 12'd2308;
    assign mem[1788] = 12'd2307;
    assign mem[1789] = 12'd2306;
    assign mem[1790] = 12'd2305;
    assign mem[1791] = 12'd2304;
    assign mem[1792] = 12'd2303;
    assign mem[1793] = 12'd2302;
    assign mem[1794] = 12'd2301;
    assign mem[1795] = 12'd2300;
    assign mem[1796] = 12'd2299;
    assign mem[1797] = 12'd2298;
    assign mem[1798] = 12'd2297;
    assign mem[1799] = 12'd2296;
    assign mem[1800] = 12'd2295;
    assign mem[1801] = 12'd2294;
    assign mem[1802] = 12'd2293;
    assign mem[1803] = 12'd2292;
    assign mem[1804] = 12'd2291;
    assign mem[1805] = 12'd2290;
    assign mem[1806] = 12'd2289;
    assign mem[1807] = 12'd2288;
    assign mem[1808] = 12'd2287;
    assign mem[1809] = 12'd2286;
    assign mem[1810] = 12'd2285;
    assign mem[1811] = 12'd2284;
    assign mem[1812] = 12'd2283;
    assign mem[1813] = 12'd2282;
    assign mem[1814] = 12'd2281;
    assign mem[1815] = 12'd2280;
    assign mem[1816] = 12'd2279;
    assign mem[1817] = 12'd2278;
    assign mem[1818] = 12'd2277;
    assign mem[1819] = 12'd2276;
    assign mem[1820] = 12'd2275;
    assign mem[1821] = 12'd2274;
    assign mem[1822] = 12'd2273;
    assign mem[1823] = 12'd2272;
    assign mem[1824] = 12'd2271;
    assign mem[1825] = 12'd2270;
    assign mem[1826] = 12'd2269;
    assign mem[1827] = 12'd2268;
    assign mem[1828] = 12'd2267;
    assign mem[1829] = 12'd2266;
    assign mem[1830] = 12'd2265;
    assign mem[1831] = 12'd2264;
    assign mem[1832] = 12'd2263;
    assign mem[1833] = 12'd2262;
    assign mem[1834] = 12'd2261;
    assign mem[1835] = 12'd2260;
    assign mem[1836] = 12'd2259;
    assign mem[1837] = 12'd2258;
    assign mem[1838] = 12'd2257;
    assign mem[1839] = 12'd2256;
    assign mem[1840] = 12'd2255;
    assign mem[1841] = 12'd2254;
    assign mem[1842] = 12'd2253;
    assign mem[1843] = 12'd2252;
    assign mem[1844] = 12'd2251;
    assign mem[1845] = 12'd2250;
    assign mem[1846] = 12'd2249;
    assign mem[1847] = 12'd2248;
    assign mem[1848] = 12'd2247;
    assign mem[1849] = 12'd2246;
    assign mem[1850] = 12'd2245;
    assign mem[1851] = 12'd2244;
    assign mem[1852] = 12'd2243;
    assign mem[1853] = 12'd2242;
    assign mem[1854] = 12'd2241;
    assign mem[1855] = 12'd2240;
    assign mem[1856] = 12'd2239;
    assign mem[1857] = 12'd2238;
    assign mem[1858] = 12'd2237;
    assign mem[1859] = 12'd2236;
    assign mem[1860] = 12'd2235;
    assign mem[1861] = 12'd2234;
    assign mem[1862] = 12'd2233;
    assign mem[1863] = 12'd2232;
    assign mem[1864] = 12'd2231;
    assign mem[1865] = 12'd2230;
    assign mem[1866] = 12'd2229;
    assign mem[1867] = 12'd2228;
    assign mem[1868] = 12'd2227;
    assign mem[1869] = 12'd2226;
    assign mem[1870] = 12'd2225;
    assign mem[1871] = 12'd2224;
    assign mem[1872] = 12'd2223;
    assign mem[1873] = 12'd2222;
    assign mem[1874] = 12'd2221;
    assign mem[1875] = 12'd2220;
    assign mem[1876] = 12'd2219;
    assign mem[1877] = 12'd2218;
    assign mem[1878] = 12'd2217;
    assign mem[1879] = 12'd2216;
    assign mem[1880] = 12'd2215;
    assign mem[1881] = 12'd2214;
    assign mem[1882] = 12'd2213;
    assign mem[1883] = 12'd2212;
    assign mem[1884] = 12'd2211;
    assign mem[1885] = 12'd2210;
    assign mem[1886] = 12'd2209;
    assign mem[1887] = 12'd2208;
    assign mem[1888] = 12'd2207;
    assign mem[1889] = 12'd2206;
    assign mem[1890] = 12'd2205;
    assign mem[1891] = 12'd2204;
    assign mem[1892] = 12'd2203;
    assign mem[1893] = 12'd2202;
    assign mem[1894] = 12'd2201;
    assign mem[1895] = 12'd2200;
    assign mem[1896] = 12'd2199;
    assign mem[1897] = 12'd2198;
    assign mem[1898] = 12'd2197;
    assign mem[1899] = 12'd2196;
    assign mem[1900] = 12'd2195;
    assign mem[1901] = 12'd2194;
    assign mem[1902] = 12'd2193;
    assign mem[1903] = 12'd2192;
    assign mem[1904] = 12'd2191;
    assign mem[1905] = 12'd2190;
    assign mem[1906] = 12'd2189;
    assign mem[1907] = 12'd2188;
    assign mem[1908] = 12'd2187;
    assign mem[1909] = 12'd2186;
    assign mem[1910] = 12'd2185;
    assign mem[1911] = 12'd2184;
    assign mem[1912] = 12'd2183;
    assign mem[1913] = 12'd2182;
    assign mem[1914] = 12'd2181;
    assign mem[1915] = 12'd2180;
    assign mem[1916] = 12'd2179;
    assign mem[1917] = 12'd2178;
    assign mem[1918] = 12'd2177;
    assign mem[1919] = 12'd2176;
    assign mem[1920] = 12'd2175;
    assign mem[1921] = 12'd2174;
    assign mem[1922] = 12'd2173;
    assign mem[1923] = 12'd2172;
    assign mem[1924] = 12'd2171;
    assign mem[1925] = 12'd2170;
    assign mem[1926] = 12'd2169;
    assign mem[1927] = 12'd2168;
    assign mem[1928] = 12'd2167;
    assign mem[1929] = 12'd2166;
    assign mem[1930] = 12'd2165;
    assign mem[1931] = 12'd2164;
    assign mem[1932] = 12'd2163;
    assign mem[1933] = 12'd2162;
    assign mem[1934] = 12'd2161;
    assign mem[1935] = 12'd2160;
    assign mem[1936] = 12'd2159;
    assign mem[1937] = 12'd2158;
    assign mem[1938] = 12'd2157;
    assign mem[1939] = 12'd2156;
    assign mem[1940] = 12'd2155;
    assign mem[1941] = 12'd2154;
    assign mem[1942] = 12'd2153;
    assign mem[1943] = 12'd2152;
    assign mem[1944] = 12'd2151;
    assign mem[1945] = 12'd2150;
    assign mem[1946] = 12'd2149;
    assign mem[1947] = 12'd2148;
    assign mem[1948] = 12'd2147;
    assign mem[1949] = 12'd2146;
    assign mem[1950] = 12'd2145;
    assign mem[1951] = 12'd2144;
    assign mem[1952] = 12'd2143;
    assign mem[1953] = 12'd2142;
    assign mem[1954] = 12'd2141;
    assign mem[1955] = 12'd2140;
    assign mem[1956] = 12'd2139;
    assign mem[1957] = 12'd2138;
    assign mem[1958] = 12'd2137;
    assign mem[1959] = 12'd2136;
    assign mem[1960] = 12'd2135;
    assign mem[1961] = 12'd2134;
    assign mem[1962] = 12'd2133;
    assign mem[1963] = 12'd2132;
    assign mem[1964] = 12'd2131;
    assign mem[1965] = 12'd2130;
    assign mem[1966] = 12'd2129;
    assign mem[1967] = 12'd2128;
    assign mem[1968] = 12'd2127;
    assign mem[1969] = 12'd2126;
    assign mem[1970] = 12'd2125;
    assign mem[1971] = 12'd2124;
    assign mem[1972] = 12'd2123;
    assign mem[1973] = 12'd2122;
    assign mem[1974] = 12'd2121;
    assign mem[1975] = 12'd2120;
    assign mem[1976] = 12'd2119;
    assign mem[1977] = 12'd2118;
    assign mem[1978] = 12'd2117;
    assign mem[1979] = 12'd2116;
    assign mem[1980] = 12'd2115;
    assign mem[1981] = 12'd2114;
    assign mem[1982] = 12'd2113;
    assign mem[1983] = 12'd2112;
    assign mem[1984] = 12'd2111;
    assign mem[1985] = 12'd2110;
    assign mem[1986] = 12'd2109;
    assign mem[1987] = 12'd2108;
    assign mem[1988] = 12'd2107;
    assign mem[1989] = 12'd2106;
    assign mem[1990] = 12'd2105;
    assign mem[1991] = 12'd2104;
    assign mem[1992] = 12'd2103;
    assign mem[1993] = 12'd2102;
    assign mem[1994] = 12'd2101;
    assign mem[1995] = 12'd2100;
    assign mem[1996] = 12'd2099;
    assign mem[1997] = 12'd2098;
    assign mem[1998] = 12'd2097;
    assign mem[1999] = 12'd2096;
    assign mem[2000] = 12'd2095;
    assign mem[2001] = 12'd2094;
    assign mem[2002] = 12'd2093;
    assign mem[2003] = 12'd2092;
    assign mem[2004] = 12'd2091;
    assign mem[2005] = 12'd2090;
    assign mem[2006] = 12'd2089;
    assign mem[2007] = 12'd2088;
    assign mem[2008] = 12'd2087;
    assign mem[2009] = 12'd2086;
    assign mem[2010] = 12'd2085;
    assign mem[2011] = 12'd2084;
    assign mem[2012] = 12'd2083;
    assign mem[2013] = 12'd2082;
    assign mem[2014] = 12'd2081;
    assign mem[2015] = 12'd2080;
    assign mem[2016] = 12'd2079;
    assign mem[2017] = 12'd2078;
    assign mem[2018] = 12'd2077;
    assign mem[2019] = 12'd2076;
    assign mem[2020] = 12'd2075;
    assign mem[2021] = 12'd2074;
    assign mem[2022] = 12'd2073;
    assign mem[2023] = 12'd2072;
    assign mem[2024] = 12'd2071;
    assign mem[2025] = 12'd2070;
    assign mem[2026] = 12'd2069;
    assign mem[2027] = 12'd2068;
    assign mem[2028] = 12'd2067;
    assign mem[2029] = 12'd2066;
    assign mem[2030] = 12'd2065;
    assign mem[2031] = 12'd2064;
    assign mem[2032] = 12'd2063;
    assign mem[2033] = 12'd2062;
    assign mem[2034] = 12'd2061;
    assign mem[2035] = 12'd2060;
    assign mem[2036] = 12'd2059;
    assign mem[2037] = 12'd2058;
    assign mem[2038] = 12'd2057;
    assign mem[2039] = 12'd2056;
    assign mem[2040] = 12'd2055;
    assign mem[2041] = 12'd2054;
    assign mem[2042] = 12'd2053;
    assign mem[2043] = 12'd2052;
    assign mem[2044] = 12'd2051;
    assign mem[2045] = 12'd2050;
    assign mem[2046] = 12'd2049;
    assign mem[2047] = 12'd2048;
    assign mem[2048] = 12'd2047;
    assign mem[2049] = 12'd2046;
    assign mem[2050] = 12'd2045;
    assign mem[2051] = 12'd2044;
    assign mem[2052] = 12'd2043;
    assign mem[2053] = 12'd2042;
    assign mem[2054] = 12'd2041;
    assign mem[2055] = 12'd2040;
    assign mem[2056] = 12'd2039;
    assign mem[2057] = 12'd2038;
    assign mem[2058] = 12'd2037;
    assign mem[2059] = 12'd2036;
    assign mem[2060] = 12'd2035;
    assign mem[2061] = 12'd2034;
    assign mem[2062] = 12'd2033;
    assign mem[2063] = 12'd2032;
    assign mem[2064] = 12'd2031;
    assign mem[2065] = 12'd2030;
    assign mem[2066] = 12'd2029;
    assign mem[2067] = 12'd2028;
    assign mem[2068] = 12'd2027;
    assign mem[2069] = 12'd2026;
    assign mem[2070] = 12'd2025;
    assign mem[2071] = 12'd2024;
    assign mem[2072] = 12'd2023;
    assign mem[2073] = 12'd2022;
    assign mem[2074] = 12'd2021;
    assign mem[2075] = 12'd2020;
    assign mem[2076] = 12'd2019;
    assign mem[2077] = 12'd2018;
    assign mem[2078] = 12'd2017;
    assign mem[2079] = 12'd2016;
    assign mem[2080] = 12'd2015;
    assign mem[2081] = 12'd2014;
    assign mem[2082] = 12'd2013;
    assign mem[2083] = 12'd2012;
    assign mem[2084] = 12'd2011;
    assign mem[2085] = 12'd2010;
    assign mem[2086] = 12'd2009;
    assign mem[2087] = 12'd2008;
    assign mem[2088] = 12'd2007;
    assign mem[2089] = 12'd2006;
    assign mem[2090] = 12'd2005;
    assign mem[2091] = 12'd2004;
    assign mem[2092] = 12'd2003;
    assign mem[2093] = 12'd2002;
    assign mem[2094] = 12'd2001;
    assign mem[2095] = 12'd2000;
    assign mem[2096] = 12'd1999;
    assign mem[2097] = 12'd1998;
    assign mem[2098] = 12'd1997;
    assign mem[2099] = 12'd1996;
    assign mem[2100] = 12'd1995;
    assign mem[2101] = 12'd1994;
    assign mem[2102] = 12'd1993;
    assign mem[2103] = 12'd1992;
    assign mem[2104] = 12'd1991;
    assign mem[2105] = 12'd1990;
    assign mem[2106] = 12'd1989;
    assign mem[2107] = 12'd1988;
    assign mem[2108] = 12'd1987;
    assign mem[2109] = 12'd1986;
    assign mem[2110] = 12'd1985;
    assign mem[2111] = 12'd1984;
    assign mem[2112] = 12'd1983;
    assign mem[2113] = 12'd1982;
    assign mem[2114] = 12'd1981;
    assign mem[2115] = 12'd1980;
    assign mem[2116] = 12'd1979;
    assign mem[2117] = 12'd1978;
    assign mem[2118] = 12'd1977;
    assign mem[2119] = 12'd1976;
    assign mem[2120] = 12'd1975;
    assign mem[2121] = 12'd1974;
    assign mem[2122] = 12'd1973;
    assign mem[2123] = 12'd1972;
    assign mem[2124] = 12'd1971;
    assign mem[2125] = 12'd1970;
    assign mem[2126] = 12'd1969;
    assign mem[2127] = 12'd1968;
    assign mem[2128] = 12'd1967;
    assign mem[2129] = 12'd1966;
    assign mem[2130] = 12'd1965;
    assign mem[2131] = 12'd1964;
    assign mem[2132] = 12'd1963;
    assign mem[2133] = 12'd1962;
    assign mem[2134] = 12'd1961;
    assign mem[2135] = 12'd1960;
    assign mem[2136] = 12'd1959;
    assign mem[2137] = 12'd1958;
    assign mem[2138] = 12'd1957;
    assign mem[2139] = 12'd1956;
    assign mem[2140] = 12'd1955;
    assign mem[2141] = 12'd1954;
    assign mem[2142] = 12'd1953;
    assign mem[2143] = 12'd1952;
    assign mem[2144] = 12'd1951;
    assign mem[2145] = 12'd1950;
    assign mem[2146] = 12'd1949;
    assign mem[2147] = 12'd1948;
    assign mem[2148] = 12'd1947;
    assign mem[2149] = 12'd1946;
    assign mem[2150] = 12'd1945;
    assign mem[2151] = 12'd1944;
    assign mem[2152] = 12'd1943;
    assign mem[2153] = 12'd1942;
    assign mem[2154] = 12'd1941;
    assign mem[2155] = 12'd1940;
    assign mem[2156] = 12'd1939;
    assign mem[2157] = 12'd1938;
    assign mem[2158] = 12'd1937;
    assign mem[2159] = 12'd1936;
    assign mem[2160] = 12'd1935;
    assign mem[2161] = 12'd1934;
    assign mem[2162] = 12'd1933;
    assign mem[2163] = 12'd1932;
    assign mem[2164] = 12'd1931;
    assign mem[2165] = 12'd1930;
    assign mem[2166] = 12'd1929;
    assign mem[2167] = 12'd1928;
    assign mem[2168] = 12'd1927;
    assign mem[2169] = 12'd1926;
    assign mem[2170] = 12'd1925;
    assign mem[2171] = 12'd1924;
    assign mem[2172] = 12'd1923;
    assign mem[2173] = 12'd1922;
    assign mem[2174] = 12'd1921;
    assign mem[2175] = 12'd1920;
    assign mem[2176] = 12'd1919;
    assign mem[2177] = 12'd1918;
    assign mem[2178] = 12'd1917;
    assign mem[2179] = 12'd1916;
    assign mem[2180] = 12'd1915;
    assign mem[2181] = 12'd1914;
    assign mem[2182] = 12'd1913;
    assign mem[2183] = 12'd1912;
    assign mem[2184] = 12'd1911;
    assign mem[2185] = 12'd1910;
    assign mem[2186] = 12'd1909;
    assign mem[2187] = 12'd1908;
    assign mem[2188] = 12'd1907;
    assign mem[2189] = 12'd1906;
    assign mem[2190] = 12'd1905;
    assign mem[2191] = 12'd1904;
    assign mem[2192] = 12'd1903;
    assign mem[2193] = 12'd1902;
    assign mem[2194] = 12'd1901;
    assign mem[2195] = 12'd1900;
    assign mem[2196] = 12'd1899;
    assign mem[2197] = 12'd1898;
    assign mem[2198] = 12'd1897;
    assign mem[2199] = 12'd1896;
    assign mem[2200] = 12'd1895;
    assign mem[2201] = 12'd1894;
    assign mem[2202] = 12'd1893;
    assign mem[2203] = 12'd1892;
    assign mem[2204] = 12'd1891;
    assign mem[2205] = 12'd1890;
    assign mem[2206] = 12'd1889;
    assign mem[2207] = 12'd1888;
    assign mem[2208] = 12'd1887;
    assign mem[2209] = 12'd1886;
    assign mem[2210] = 12'd1885;
    assign mem[2211] = 12'd1884;
    assign mem[2212] = 12'd1883;
    assign mem[2213] = 12'd1882;
    assign mem[2214] = 12'd1881;
    assign mem[2215] = 12'd1880;
    assign mem[2216] = 12'd1879;
    assign mem[2217] = 12'd1878;
    assign mem[2218] = 12'd1877;
    assign mem[2219] = 12'd1876;
    assign mem[2220] = 12'd1875;
    assign mem[2221] = 12'd1874;
    assign mem[2222] = 12'd1873;
    assign mem[2223] = 12'd1872;
    assign mem[2224] = 12'd1871;
    assign mem[2225] = 12'd1870;
    assign mem[2226] = 12'd1869;
    assign mem[2227] = 12'd1868;
    assign mem[2228] = 12'd1867;
    assign mem[2229] = 12'd1866;
    assign mem[2230] = 12'd1865;
    assign mem[2231] = 12'd1864;
    assign mem[2232] = 12'd1863;
    assign mem[2233] = 12'd1862;
    assign mem[2234] = 12'd1861;
    assign mem[2235] = 12'd1860;
    assign mem[2236] = 12'd1859;
    assign mem[2237] = 12'd1858;
    assign mem[2238] = 12'd1857;
    assign mem[2239] = 12'd1856;
    assign mem[2240] = 12'd1855;
    assign mem[2241] = 12'd1854;
    assign mem[2242] = 12'd1853;
    assign mem[2243] = 12'd1852;
    assign mem[2244] = 12'd1851;
    assign mem[2245] = 12'd1850;
    assign mem[2246] = 12'd1849;
    assign mem[2247] = 12'd1848;
    assign mem[2248] = 12'd1847;
    assign mem[2249] = 12'd1846;
    assign mem[2250] = 12'd1845;
    assign mem[2251] = 12'd1844;
    assign mem[2252] = 12'd1843;
    assign mem[2253] = 12'd1842;
    assign mem[2254] = 12'd1841;
    assign mem[2255] = 12'd1840;
    assign mem[2256] = 12'd1839;
    assign mem[2257] = 12'd1838;
    assign mem[2258] = 12'd1837;
    assign mem[2259] = 12'd1836;
    assign mem[2260] = 12'd1835;
    assign mem[2261] = 12'd1834;
    assign mem[2262] = 12'd1833;
    assign mem[2263] = 12'd1832;
    assign mem[2264] = 12'd1831;
    assign mem[2265] = 12'd1830;
    assign mem[2266] = 12'd1829;
    assign mem[2267] = 12'd1828;
    assign mem[2268] = 12'd1827;
    assign mem[2269] = 12'd1826;
    assign mem[2270] = 12'd1825;
    assign mem[2271] = 12'd1824;
    assign mem[2272] = 12'd1823;
    assign mem[2273] = 12'd1822;
    assign mem[2274] = 12'd1821;
    assign mem[2275] = 12'd1820;
    assign mem[2276] = 12'd1819;
    assign mem[2277] = 12'd1818;
    assign mem[2278] = 12'd1817;
    assign mem[2279] = 12'd1816;
    assign mem[2280] = 12'd1815;
    assign mem[2281] = 12'd1814;
    assign mem[2282] = 12'd1813;
    assign mem[2283] = 12'd1812;
    assign mem[2284] = 12'd1811;
    assign mem[2285] = 12'd1810;
    assign mem[2286] = 12'd1809;
    assign mem[2287] = 12'd1808;
    assign mem[2288] = 12'd1807;
    assign mem[2289] = 12'd1806;
    assign mem[2290] = 12'd1805;
    assign mem[2291] = 12'd1804;
    assign mem[2292] = 12'd1803;
    assign mem[2293] = 12'd1802;
    assign mem[2294] = 12'd1801;
    assign mem[2295] = 12'd1800;
    assign mem[2296] = 12'd1799;
    assign mem[2297] = 12'd1798;
    assign mem[2298] = 12'd1797;
    assign mem[2299] = 12'd1796;
    assign mem[2300] = 12'd1795;
    assign mem[2301] = 12'd1794;
    assign mem[2302] = 12'd1793;
    assign mem[2303] = 12'd1792;
    assign mem[2304] = 12'd1791;
    assign mem[2305] = 12'd1790;
    assign mem[2306] = 12'd1789;
    assign mem[2307] = 12'd1788;
    assign mem[2308] = 12'd1787;
    assign mem[2309] = 12'd1786;
    assign mem[2310] = 12'd1785;
    assign mem[2311] = 12'd1784;
    assign mem[2312] = 12'd1783;
    assign mem[2313] = 12'd1782;
    assign mem[2314] = 12'd1781;
    assign mem[2315] = 12'd1780;
    assign mem[2316] = 12'd1779;
    assign mem[2317] = 12'd1778;
    assign mem[2318] = 12'd1777;
    assign mem[2319] = 12'd1776;
    assign mem[2320] = 12'd1775;
    assign mem[2321] = 12'd1774;
    assign mem[2322] = 12'd1773;
    assign mem[2323] = 12'd1772;
    assign mem[2324] = 12'd1771;
    assign mem[2325] = 12'd1770;
    assign mem[2326] = 12'd1769;
    assign mem[2327] = 12'd1768;
    assign mem[2328] = 12'd1767;
    assign mem[2329] = 12'd1766;
    assign mem[2330] = 12'd1765;
    assign mem[2331] = 12'd1764;
    assign mem[2332] = 12'd1763;
    assign mem[2333] = 12'd1762;
    assign mem[2334] = 12'd1761;
    assign mem[2335] = 12'd1760;
    assign mem[2336] = 12'd1759;
    assign mem[2337] = 12'd1758;
    assign mem[2338] = 12'd1757;
    assign mem[2339] = 12'd1756;
    assign mem[2340] = 12'd1755;
    assign mem[2341] = 12'd1754;
    assign mem[2342] = 12'd1753;
    assign mem[2343] = 12'd1752;
    assign mem[2344] = 12'd1751;
    assign mem[2345] = 12'd1750;
    assign mem[2346] = 12'd1749;
    assign mem[2347] = 12'd1748;
    assign mem[2348] = 12'd1747;
    assign mem[2349] = 12'd1746;
    assign mem[2350] = 12'd1745;
    assign mem[2351] = 12'd1744;
    assign mem[2352] = 12'd1743;
    assign mem[2353] = 12'd1742;
    assign mem[2354] = 12'd1741;
    assign mem[2355] = 12'd1740;
    assign mem[2356] = 12'd1739;
    assign mem[2357] = 12'd1738;
    assign mem[2358] = 12'd1737;
    assign mem[2359] = 12'd1736;
    assign mem[2360] = 12'd1735;
    assign mem[2361] = 12'd1734;
    assign mem[2362] = 12'd1733;
    assign mem[2363] = 12'd1732;
    assign mem[2364] = 12'd1731;
    assign mem[2365] = 12'd1730;
    assign mem[2366] = 12'd1729;
    assign mem[2367] = 12'd1728;
    assign mem[2368] = 12'd1727;
    assign mem[2369] = 12'd1726;
    assign mem[2370] = 12'd1725;
    assign mem[2371] = 12'd1724;
    assign mem[2372] = 12'd1723;
    assign mem[2373] = 12'd1722;
    assign mem[2374] = 12'd1721;
    assign mem[2375] = 12'd1720;
    assign mem[2376] = 12'd1719;
    assign mem[2377] = 12'd1718;
    assign mem[2378] = 12'd1717;
    assign mem[2379] = 12'd1716;
    assign mem[2380] = 12'd1715;
    assign mem[2381] = 12'd1714;
    assign mem[2382] = 12'd1713;
    assign mem[2383] = 12'd1712;
    assign mem[2384] = 12'd1711;
    assign mem[2385] = 12'd1710;
    assign mem[2386] = 12'd1709;
    assign mem[2387] = 12'd1708;
    assign mem[2388] = 12'd1707;
    assign mem[2389] = 12'd1706;
    assign mem[2390] = 12'd1705;
    assign mem[2391] = 12'd1704;
    assign mem[2392] = 12'd1703;
    assign mem[2393] = 12'd1702;
    assign mem[2394] = 12'd1701;
    assign mem[2395] = 12'd1700;
    assign mem[2396] = 12'd1699;
    assign mem[2397] = 12'd1698;
    assign mem[2398] = 12'd1697;
    assign mem[2399] = 12'd1696;
    assign mem[2400] = 12'd1695;
    assign mem[2401] = 12'd1694;
    assign mem[2402] = 12'd1693;
    assign mem[2403] = 12'd1692;
    assign mem[2404] = 12'd1691;
    assign mem[2405] = 12'd1690;
    assign mem[2406] = 12'd1689;
    assign mem[2407] = 12'd1688;
    assign mem[2408] = 12'd1687;
    assign mem[2409] = 12'd1686;
    assign mem[2410] = 12'd1685;
    assign mem[2411] = 12'd1684;
    assign mem[2412] = 12'd1683;
    assign mem[2413] = 12'd1682;
    assign mem[2414] = 12'd1681;
    assign mem[2415] = 12'd1680;
    assign mem[2416] = 12'd1679;
    assign mem[2417] = 12'd1678;
    assign mem[2418] = 12'd1677;
    assign mem[2419] = 12'd1676;
    assign mem[2420] = 12'd1675;
    assign mem[2421] = 12'd1674;
    assign mem[2422] = 12'd1673;
    assign mem[2423] = 12'd1672;
    assign mem[2424] = 12'd1671;
    assign mem[2425] = 12'd1670;
    assign mem[2426] = 12'd1669;
    assign mem[2427] = 12'd1668;
    assign mem[2428] = 12'd1667;
    assign mem[2429] = 12'd1666;
    assign mem[2430] = 12'd1665;
    assign mem[2431] = 12'd1664;
    assign mem[2432] = 12'd1663;
    assign mem[2433] = 12'd1662;
    assign mem[2434] = 12'd1661;
    assign mem[2435] = 12'd1660;
    assign mem[2436] = 12'd1659;
    assign mem[2437] = 12'd1658;
    assign mem[2438] = 12'd1657;
    assign mem[2439] = 12'd1656;
    assign mem[2440] = 12'd1655;
    assign mem[2441] = 12'd1654;
    assign mem[2442] = 12'd1653;
    assign mem[2443] = 12'd1652;
    assign mem[2444] = 12'd1651;
    assign mem[2445] = 12'd1650;
    assign mem[2446] = 12'd1649;
    assign mem[2447] = 12'd1648;
    assign mem[2448] = 12'd1647;
    assign mem[2449] = 12'd1646;
    assign mem[2450] = 12'd1645;
    assign mem[2451] = 12'd1644;
    assign mem[2452] = 12'd1643;
    assign mem[2453] = 12'd1642;
    assign mem[2454] = 12'd1641;
    assign mem[2455] = 12'd1640;
    assign mem[2456] = 12'd1639;
    assign mem[2457] = 12'd1638;
    assign mem[2458] = 12'd1637;
    assign mem[2459] = 12'd1636;
    assign mem[2460] = 12'd1635;
    assign mem[2461] = 12'd1634;
    assign mem[2462] = 12'd1633;
    assign mem[2463] = 12'd1632;
    assign mem[2464] = 12'd1631;
    assign mem[2465] = 12'd1630;
    assign mem[2466] = 12'd1629;
    assign mem[2467] = 12'd1628;
    assign mem[2468] = 12'd1627;
    assign mem[2469] = 12'd1626;
    assign mem[2470] = 12'd1625;
    assign mem[2471] = 12'd1624;
    assign mem[2472] = 12'd1623;
    assign mem[2473] = 12'd1622;
    assign mem[2474] = 12'd1621;
    assign mem[2475] = 12'd1620;
    assign mem[2476] = 12'd1619;
    assign mem[2477] = 12'd1618;
    assign mem[2478] = 12'd1617;
    assign mem[2479] = 12'd1616;
    assign mem[2480] = 12'd1615;
    assign mem[2481] = 12'd1614;
    assign mem[2482] = 12'd1613;
    assign mem[2483] = 12'd1612;
    assign mem[2484] = 12'd1611;
    assign mem[2485] = 12'd1610;
    assign mem[2486] = 12'd1609;
    assign mem[2487] = 12'd1608;
    assign mem[2488] = 12'd1607;
    assign mem[2489] = 12'd1606;
    assign mem[2490] = 12'd1605;
    assign mem[2491] = 12'd1604;
    assign mem[2492] = 12'd1603;
    assign mem[2493] = 12'd1602;
    assign mem[2494] = 12'd1601;
    assign mem[2495] = 12'd1600;
    assign mem[2496] = 12'd1599;
    assign mem[2497] = 12'd1598;
    assign mem[2498] = 12'd1597;
    assign mem[2499] = 12'd1596;
    assign mem[2500] = 12'd1595;
    assign mem[2501] = 12'd1594;
    assign mem[2502] = 12'd1593;
    assign mem[2503] = 12'd1592;
    assign mem[2504] = 12'd1591;
    assign mem[2505] = 12'd1590;
    assign mem[2506] = 12'd1589;
    assign mem[2507] = 12'd1588;
    assign mem[2508] = 12'd1587;
    assign mem[2509] = 12'd1586;
    assign mem[2510] = 12'd1585;
    assign mem[2511] = 12'd1584;
    assign mem[2512] = 12'd1583;
    assign mem[2513] = 12'd1582;
    assign mem[2514] = 12'd1581;
    assign mem[2515] = 12'd1580;
    assign mem[2516] = 12'd1579;
    assign mem[2517] = 12'd1578;
    assign mem[2518] = 12'd1577;
    assign mem[2519] = 12'd1576;
    assign mem[2520] = 12'd1575;
    assign mem[2521] = 12'd1574;
    assign mem[2522] = 12'd1573;
    assign mem[2523] = 12'd1572;
    assign mem[2524] = 12'd1571;
    assign mem[2525] = 12'd1570;
    assign mem[2526] = 12'd1569;
    assign mem[2527] = 12'd1568;
    assign mem[2528] = 12'd1567;
    assign mem[2529] = 12'd1566;
    assign mem[2530] = 12'd1565;
    assign mem[2531] = 12'd1564;
    assign mem[2532] = 12'd1563;
    assign mem[2533] = 12'd1562;
    assign mem[2534] = 12'd1561;
    assign mem[2535] = 12'd1560;
    assign mem[2536] = 12'd1559;
    assign mem[2537] = 12'd1558;
    assign mem[2538] = 12'd1557;
    assign mem[2539] = 12'd1556;
    assign mem[2540] = 12'd1555;
    assign mem[2541] = 12'd1554;
    assign mem[2542] = 12'd1553;
    assign mem[2543] = 12'd1552;
    assign mem[2544] = 12'd1551;
    assign mem[2545] = 12'd1550;
    assign mem[2546] = 12'd1549;
    assign mem[2547] = 12'd1548;
    assign mem[2548] = 12'd1547;
    assign mem[2549] = 12'd1546;
    assign mem[2550] = 12'd1545;
    assign mem[2551] = 12'd1544;
    assign mem[2552] = 12'd1543;
    assign mem[2553] = 12'd1542;
    assign mem[2554] = 12'd1541;
    assign mem[2555] = 12'd1540;
    assign mem[2556] = 12'd1539;
    assign mem[2557] = 12'd1538;
    assign mem[2558] = 12'd1537;
    assign mem[2559] = 12'd1536;
    assign mem[2560] = 12'd1535;
    assign mem[2561] = 12'd1534;
    assign mem[2562] = 12'd1533;
    assign mem[2563] = 12'd1532;
    assign mem[2564] = 12'd1531;
    assign mem[2565] = 12'd1530;
    assign mem[2566] = 12'd1529;
    assign mem[2567] = 12'd1528;
    assign mem[2568] = 12'd1527;
    assign mem[2569] = 12'd1526;
    assign mem[2570] = 12'd1525;
    assign mem[2571] = 12'd1524;
    assign mem[2572] = 12'd1523;
    assign mem[2573] = 12'd1522;
    assign mem[2574] = 12'd1521;
    assign mem[2575] = 12'd1520;
    assign mem[2576] = 12'd1519;
    assign mem[2577] = 12'd1518;
    assign mem[2578] = 12'd1517;
    assign mem[2579] = 12'd1516;
    assign mem[2580] = 12'd1515;
    assign mem[2581] = 12'd1514;
    assign mem[2582] = 12'd1513;
    assign mem[2583] = 12'd1512;
    assign mem[2584] = 12'd1511;
    assign mem[2585] = 12'd1510;
    assign mem[2586] = 12'd1509;
    assign mem[2587] = 12'd1508;
    assign mem[2588] = 12'd1507;
    assign mem[2589] = 12'd1506;
    assign mem[2590] = 12'd1505;
    assign mem[2591] = 12'd1504;
    assign mem[2592] = 12'd1503;
    assign mem[2593] = 12'd1502;
    assign mem[2594] = 12'd1501;
    assign mem[2595] = 12'd1500;
    assign mem[2596] = 12'd1499;
    assign mem[2597] = 12'd1498;
    assign mem[2598] = 12'd1497;
    assign mem[2599] = 12'd1496;
    assign mem[2600] = 12'd1495;
    assign mem[2601] = 12'd1494;
    assign mem[2602] = 12'd1493;
    assign mem[2603] = 12'd1492;
    assign mem[2604] = 12'd1491;
    assign mem[2605] = 12'd1490;
    assign mem[2606] = 12'd1489;
    assign mem[2607] = 12'd1488;
    assign mem[2608] = 12'd1487;
    assign mem[2609] = 12'd1486;
    assign mem[2610] = 12'd1485;
    assign mem[2611] = 12'd1484;
    assign mem[2612] = 12'd1483;
    assign mem[2613] = 12'd1482;
    assign mem[2614] = 12'd1481;
    assign mem[2615] = 12'd1480;
    assign mem[2616] = 12'd1479;
    assign mem[2617] = 12'd1478;
    assign mem[2618] = 12'd1477;
    assign mem[2619] = 12'd1476;
    assign mem[2620] = 12'd1475;
    assign mem[2621] = 12'd1474;
    assign mem[2622] = 12'd1473;
    assign mem[2623] = 12'd1472;
    assign mem[2624] = 12'd1471;
    assign mem[2625] = 12'd1470;
    assign mem[2626] = 12'd1469;
    assign mem[2627] = 12'd1468;
    assign mem[2628] = 12'd1467;
    assign mem[2629] = 12'd1466;
    assign mem[2630] = 12'd1465;
    assign mem[2631] = 12'd1464;
    assign mem[2632] = 12'd1463;
    assign mem[2633] = 12'd1462;
    assign mem[2634] = 12'd1461;
    assign mem[2635] = 12'd1460;
    assign mem[2636] = 12'd1459;
    assign mem[2637] = 12'd1458;
    assign mem[2638] = 12'd1457;
    assign mem[2639] = 12'd1456;
    assign mem[2640] = 12'd1455;
    assign mem[2641] = 12'd1454;
    assign mem[2642] = 12'd1453;
    assign mem[2643] = 12'd1452;
    assign mem[2644] = 12'd1451;
    assign mem[2645] = 12'd1450;
    assign mem[2646] = 12'd1449;
    assign mem[2647] = 12'd1448;
    assign mem[2648] = 12'd1447;
    assign mem[2649] = 12'd1446;
    assign mem[2650] = 12'd1445;
    assign mem[2651] = 12'd1444;
    assign mem[2652] = 12'd1443;
    assign mem[2653] = 12'd1442;
    assign mem[2654] = 12'd1441;
    assign mem[2655] = 12'd1440;
    assign mem[2656] = 12'd1439;
    assign mem[2657] = 12'd1438;
    assign mem[2658] = 12'd1437;
    assign mem[2659] = 12'd1436;
    assign mem[2660] = 12'd1435;
    assign mem[2661] = 12'd1434;
    assign mem[2662] = 12'd1433;
    assign mem[2663] = 12'd1432;
    assign mem[2664] = 12'd1431;
    assign mem[2665] = 12'd1430;
    assign mem[2666] = 12'd1429;
    assign mem[2667] = 12'd1428;
    assign mem[2668] = 12'd1427;
    assign mem[2669] = 12'd1426;
    assign mem[2670] = 12'd1425;
    assign mem[2671] = 12'd1424;
    assign mem[2672] = 12'd1423;
    assign mem[2673] = 12'd1422;
    assign mem[2674] = 12'd1421;
    assign mem[2675] = 12'd1420;
    assign mem[2676] = 12'd1419;
    assign mem[2677] = 12'd1418;
    assign mem[2678] = 12'd1417;
    assign mem[2679] = 12'd1416;
    assign mem[2680] = 12'd1415;
    assign mem[2681] = 12'd1414;
    assign mem[2682] = 12'd1413;
    assign mem[2683] = 12'd1412;
    assign mem[2684] = 12'd1411;
    assign mem[2685] = 12'd1410;
    assign mem[2686] = 12'd1409;
    assign mem[2687] = 12'd1408;
    assign mem[2688] = 12'd1407;
    assign mem[2689] = 12'd1406;
    assign mem[2690] = 12'd1405;
    assign mem[2691] = 12'd1404;
    assign mem[2692] = 12'd1403;
    assign mem[2693] = 12'd1402;
    assign mem[2694] = 12'd1401;
    assign mem[2695] = 12'd1400;
    assign mem[2696] = 12'd1399;
    assign mem[2697] = 12'd1398;
    assign mem[2698] = 12'd1397;
    assign mem[2699] = 12'd1396;
    assign mem[2700] = 12'd1395;
    assign mem[2701] = 12'd1394;
    assign mem[2702] = 12'd1393;
    assign mem[2703] = 12'd1392;
    assign mem[2704] = 12'd1391;
    assign mem[2705] = 12'd1390;
    assign mem[2706] = 12'd1389;
    assign mem[2707] = 12'd1388;
    assign mem[2708] = 12'd1387;
    assign mem[2709] = 12'd1386;
    assign mem[2710] = 12'd1385;
    assign mem[2711] = 12'd1384;
    assign mem[2712] = 12'd1383;
    assign mem[2713] = 12'd1382;
    assign mem[2714] = 12'd1381;
    assign mem[2715] = 12'd1380;
    assign mem[2716] = 12'd1379;
    assign mem[2717] = 12'd1378;
    assign mem[2718] = 12'd1377;
    assign mem[2719] = 12'd1376;
    assign mem[2720] = 12'd1375;
    assign mem[2721] = 12'd1374;
    assign mem[2722] = 12'd1373;
    assign mem[2723] = 12'd1372;
    assign mem[2724] = 12'd1371;
    assign mem[2725] = 12'd1370;
    assign mem[2726] = 12'd1369;
    assign mem[2727] = 12'd1368;
    assign mem[2728] = 12'd1367;
    assign mem[2729] = 12'd1366;
    assign mem[2730] = 12'd1365;
    assign mem[2731] = 12'd1364;
    assign mem[2732] = 12'd1363;
    assign mem[2733] = 12'd1362;
    assign mem[2734] = 12'd1361;
    assign mem[2735] = 12'd1360;
    assign mem[2736] = 12'd1359;
    assign mem[2737] = 12'd1358;
    assign mem[2738] = 12'd1357;
    assign mem[2739] = 12'd1356;
    assign mem[2740] = 12'd1355;
    assign mem[2741] = 12'd1354;
    assign mem[2742] = 12'd1353;
    assign mem[2743] = 12'd1352;
    assign mem[2744] = 12'd1351;
    assign mem[2745] = 12'd1350;
    assign mem[2746] = 12'd1349;
    assign mem[2747] = 12'd1348;
    assign mem[2748] = 12'd1347;
    assign mem[2749] = 12'd1346;
    assign mem[2750] = 12'd1345;
    assign mem[2751] = 12'd1344;
    assign mem[2752] = 12'd1343;
    assign mem[2753] = 12'd1342;
    assign mem[2754] = 12'd1341;
    assign mem[2755] = 12'd1340;
    assign mem[2756] = 12'd1339;
    assign mem[2757] = 12'd1338;
    assign mem[2758] = 12'd1337;
    assign mem[2759] = 12'd1336;
    assign mem[2760] = 12'd1335;
    assign mem[2761] = 12'd1334;
    assign mem[2762] = 12'd1333;
    assign mem[2763] = 12'd1332;
    assign mem[2764] = 12'd1331;
    assign mem[2765] = 12'd1330;
    assign mem[2766] = 12'd1329;
    assign mem[2767] = 12'd1328;
    assign mem[2768] = 12'd1327;
    assign mem[2769] = 12'd1326;
    assign mem[2770] = 12'd1325;
    assign mem[2771] = 12'd1324;
    assign mem[2772] = 12'd1323;
    assign mem[2773] = 12'd1322;
    assign mem[2774] = 12'd1321;
    assign mem[2775] = 12'd1320;
    assign mem[2776] = 12'd1319;
    assign mem[2777] = 12'd1318;
    assign mem[2778] = 12'd1317;
    assign mem[2779] = 12'd1316;
    assign mem[2780] = 12'd1315;
    assign mem[2781] = 12'd1314;
    assign mem[2782] = 12'd1313;
    assign mem[2783] = 12'd1312;
    assign mem[2784] = 12'd1311;
    assign mem[2785] = 12'd1310;
    assign mem[2786] = 12'd1309;
    assign mem[2787] = 12'd1308;
    assign mem[2788] = 12'd1307;
    assign mem[2789] = 12'd1306;
    assign mem[2790] = 12'd1305;
    assign mem[2791] = 12'd1304;
    assign mem[2792] = 12'd1303;
    assign mem[2793] = 12'd1302;
    assign mem[2794] = 12'd1301;
    assign mem[2795] = 12'd1300;
    assign mem[2796] = 12'd1299;
    assign mem[2797] = 12'd1298;
    assign mem[2798] = 12'd1297;
    assign mem[2799] = 12'd1296;
    assign mem[2800] = 12'd1295;
    assign mem[2801] = 12'd1294;
    assign mem[2802] = 12'd1293;
    assign mem[2803] = 12'd1292;
    assign mem[2804] = 12'd1291;
    assign mem[2805] = 12'd1290;
    assign mem[2806] = 12'd1289;
    assign mem[2807] = 12'd1288;
    assign mem[2808] = 12'd1287;
    assign mem[2809] = 12'd1286;
    assign mem[2810] = 12'd1285;
    assign mem[2811] = 12'd1284;
    assign mem[2812] = 12'd1283;
    assign mem[2813] = 12'd1282;
    assign mem[2814] = 12'd1281;
    assign mem[2815] = 12'd1280;
    assign mem[2816] = 12'd1279;
    assign mem[2817] = 12'd1278;
    assign mem[2818] = 12'd1277;
    assign mem[2819] = 12'd1276;
    assign mem[2820] = 12'd1275;
    assign mem[2821] = 12'd1274;
    assign mem[2822] = 12'd1273;
    assign mem[2823] = 12'd1272;
    assign mem[2824] = 12'd1271;
    assign mem[2825] = 12'd1270;
    assign mem[2826] = 12'd1269;
    assign mem[2827] = 12'd1268;
    assign mem[2828] = 12'd1267;
    assign mem[2829] = 12'd1266;
    assign mem[2830] = 12'd1265;
    assign mem[2831] = 12'd1264;
    assign mem[2832] = 12'd1263;
    assign mem[2833] = 12'd1262;
    assign mem[2834] = 12'd1261;
    assign mem[2835] = 12'd1260;
    assign mem[2836] = 12'd1259;
    assign mem[2837] = 12'd1258;
    assign mem[2838] = 12'd1257;
    assign mem[2839] = 12'd1256;
    assign mem[2840] = 12'd1255;
    assign mem[2841] = 12'd1254;
    assign mem[2842] = 12'd1253;
    assign mem[2843] = 12'd1252;
    assign mem[2844] = 12'd1251;
    assign mem[2845] = 12'd1250;
    assign mem[2846] = 12'd1249;
    assign mem[2847] = 12'd1248;
    assign mem[2848] = 12'd1247;
    assign mem[2849] = 12'd1246;
    assign mem[2850] = 12'd1245;
    assign mem[2851] = 12'd1244;
    assign mem[2852] = 12'd1243;
    assign mem[2853] = 12'd1242;
    assign mem[2854] = 12'd1241;
    assign mem[2855] = 12'd1240;
    assign mem[2856] = 12'd1239;
    assign mem[2857] = 12'd1238;
    assign mem[2858] = 12'd1237;
    assign mem[2859] = 12'd1236;
    assign mem[2860] = 12'd1235;
    assign mem[2861] = 12'd1234;
    assign mem[2862] = 12'd1233;
    assign mem[2863] = 12'd1232;
    assign mem[2864] = 12'd1231;
    assign mem[2865] = 12'd1230;
    assign mem[2866] = 12'd1229;
    assign mem[2867] = 12'd1228;
    assign mem[2868] = 12'd1227;
    assign mem[2869] = 12'd1226;
    assign mem[2870] = 12'd1225;
    assign mem[2871] = 12'd1224;
    assign mem[2872] = 12'd1223;
    assign mem[2873] = 12'd1222;
    assign mem[2874] = 12'd1221;
    assign mem[2875] = 12'd1220;
    assign mem[2876] = 12'd1219;
    assign mem[2877] = 12'd1218;
    assign mem[2878] = 12'd1217;
    assign mem[2879] = 12'd1216;
    assign mem[2880] = 12'd1215;
    assign mem[2881] = 12'd1214;
    assign mem[2882] = 12'd1213;
    assign mem[2883] = 12'd1212;
    assign mem[2884] = 12'd1211;
    assign mem[2885] = 12'd1210;
    assign mem[2886] = 12'd1209;
    assign mem[2887] = 12'd1208;
    assign mem[2888] = 12'd1207;
    assign mem[2889] = 12'd1206;
    assign mem[2890] = 12'd1205;
    assign mem[2891] = 12'd1204;
    assign mem[2892] = 12'd1203;
    assign mem[2893] = 12'd1202;
    assign mem[2894] = 12'd1201;
    assign mem[2895] = 12'd1200;
    assign mem[2896] = 12'd1199;
    assign mem[2897] = 12'd1198;
    assign mem[2898] = 12'd1197;
    assign mem[2899] = 12'd1196;
    assign mem[2900] = 12'd1195;
    assign mem[2901] = 12'd1194;
    assign mem[2902] = 12'd1193;
    assign mem[2903] = 12'd1192;
    assign mem[2904] = 12'd1191;
    assign mem[2905] = 12'd1190;
    assign mem[2906] = 12'd1189;
    assign mem[2907] = 12'd1188;
    assign mem[2908] = 12'd1187;
    assign mem[2909] = 12'd1186;
    assign mem[2910] = 12'd1185;
    assign mem[2911] = 12'd1184;
    assign mem[2912] = 12'd1183;
    assign mem[2913] = 12'd1182;
    assign mem[2914] = 12'd1181;
    assign mem[2915] = 12'd1180;
    assign mem[2916] = 12'd1179;
    assign mem[2917] = 12'd1178;
    assign mem[2918] = 12'd1177;
    assign mem[2919] = 12'd1176;
    assign mem[2920] = 12'd1175;
    assign mem[2921] = 12'd1174;
    assign mem[2922] = 12'd1173;
    assign mem[2923] = 12'd1172;
    assign mem[2924] = 12'd1171;
    assign mem[2925] = 12'd1170;
    assign mem[2926] = 12'd1169;
    assign mem[2927] = 12'd1168;
    assign mem[2928] = 12'd1167;
    assign mem[2929] = 12'd1166;
    assign mem[2930] = 12'd1165;
    assign mem[2931] = 12'd1164;
    assign mem[2932] = 12'd1163;
    assign mem[2933] = 12'd1162;
    assign mem[2934] = 12'd1161;
    assign mem[2935] = 12'd1160;
    assign mem[2936] = 12'd1159;
    assign mem[2937] = 12'd1158;
    assign mem[2938] = 12'd1157;
    assign mem[2939] = 12'd1156;
    assign mem[2940] = 12'd1155;
    assign mem[2941] = 12'd1154;
    assign mem[2942] = 12'd1153;
    assign mem[2943] = 12'd1152;
    assign mem[2944] = 12'd1151;
    assign mem[2945] = 12'd1150;
    assign mem[2946] = 12'd1149;
    assign mem[2947] = 12'd1148;
    assign mem[2948] = 12'd1147;
    assign mem[2949] = 12'd1146;
    assign mem[2950] = 12'd1145;
    assign mem[2951] = 12'd1144;
    assign mem[2952] = 12'd1143;
    assign mem[2953] = 12'd1142;
    assign mem[2954] = 12'd1141;
    assign mem[2955] = 12'd1140;
    assign mem[2956] = 12'd1139;
    assign mem[2957] = 12'd1138;
    assign mem[2958] = 12'd1137;
    assign mem[2959] = 12'd1136;
    assign mem[2960] = 12'd1135;
    assign mem[2961] = 12'd1134;
    assign mem[2962] = 12'd1133;
    assign mem[2963] = 12'd1132;
    assign mem[2964] = 12'd1131;
    assign mem[2965] = 12'd1130;
    assign mem[2966] = 12'd1129;
    assign mem[2967] = 12'd1128;
    assign mem[2968] = 12'd1127;
    assign mem[2969] = 12'd1126;
    assign mem[2970] = 12'd1125;
    assign mem[2971] = 12'd1124;
    assign mem[2972] = 12'd1123;
    assign mem[2973] = 12'd1122;
    assign mem[2974] = 12'd1121;
    assign mem[2975] = 12'd1120;
    assign mem[2976] = 12'd1119;
    assign mem[2977] = 12'd1118;
    assign mem[2978] = 12'd1117;
    assign mem[2979] = 12'd1116;
    assign mem[2980] = 12'd1115;
    assign mem[2981] = 12'd1114;
    assign mem[2982] = 12'd1113;
    assign mem[2983] = 12'd1112;
    assign mem[2984] = 12'd1111;
    assign mem[2985] = 12'd1110;
    assign mem[2986] = 12'd1109;
    assign mem[2987] = 12'd1108;
    assign mem[2988] = 12'd1107;
    assign mem[2989] = 12'd1106;
    assign mem[2990] = 12'd1105;
    assign mem[2991] = 12'd1104;
    assign mem[2992] = 12'd1103;
    assign mem[2993] = 12'd1102;
    assign mem[2994] = 12'd1101;
    assign mem[2995] = 12'd1100;
    assign mem[2996] = 12'd1099;
    assign mem[2997] = 12'd1098;
    assign mem[2998] = 12'd1097;
    assign mem[2999] = 12'd1096;
    assign mem[3000] = 12'd1095;
    assign mem[3001] = 12'd1094;
    assign mem[3002] = 12'd1093;
    assign mem[3003] = 12'd1092;
    assign mem[3004] = 12'd1091;
    assign mem[3005] = 12'd1090;
    assign mem[3006] = 12'd1089;
    assign mem[3007] = 12'd1088;
    assign mem[3008] = 12'd1087;
    assign mem[3009] = 12'd1086;
    assign mem[3010] = 12'd1085;
    assign mem[3011] = 12'd1084;
    assign mem[3012] = 12'd1083;
    assign mem[3013] = 12'd1082;
    assign mem[3014] = 12'd1081;
    assign mem[3015] = 12'd1080;
    assign mem[3016] = 12'd1079;
    assign mem[3017] = 12'd1078;
    assign mem[3018] = 12'd1077;
    assign mem[3019] = 12'd1076;
    assign mem[3020] = 12'd1075;
    assign mem[3021] = 12'd1074;
    assign mem[3022] = 12'd1073;
    assign mem[3023] = 12'd1072;
    assign mem[3024] = 12'd1071;
    assign mem[3025] = 12'd1070;
    assign mem[3026] = 12'd1069;
    assign mem[3027] = 12'd1068;
    assign mem[3028] = 12'd1067;
    assign mem[3029] = 12'd1066;
    assign mem[3030] = 12'd1065;
    assign mem[3031] = 12'd1064;
    assign mem[3032] = 12'd1063;
    assign mem[3033] = 12'd1062;
    assign mem[3034] = 12'd1061;
    assign mem[3035] = 12'd1060;
    assign mem[3036] = 12'd1059;
    assign mem[3037] = 12'd1058;
    assign mem[3038] = 12'd1057;
    assign mem[3039] = 12'd1056;
    assign mem[3040] = 12'd1055;
    assign mem[3041] = 12'd1054;
    assign mem[3042] = 12'd1053;
    assign mem[3043] = 12'd1052;
    assign mem[3044] = 12'd1051;
    assign mem[3045] = 12'd1050;
    assign mem[3046] = 12'd1049;
    assign mem[3047] = 12'd1048;
    assign mem[3048] = 12'd1047;
    assign mem[3049] = 12'd1046;
    assign mem[3050] = 12'd1045;
    assign mem[3051] = 12'd1044;
    assign mem[3052] = 12'd1043;
    assign mem[3053] = 12'd1042;
    assign mem[3054] = 12'd1041;
    assign mem[3055] = 12'd1040;
    assign mem[3056] = 12'd1039;
    assign mem[3057] = 12'd1038;
    assign mem[3058] = 12'd1037;
    assign mem[3059] = 12'd1036;
    assign mem[3060] = 12'd1035;
    assign mem[3061] = 12'd1034;
    assign mem[3062] = 12'd1033;
    assign mem[3063] = 12'd1032;
    assign mem[3064] = 12'd1031;
    assign mem[3065] = 12'd1030;
    assign mem[3066] = 12'd1029;
    assign mem[3067] = 12'd1028;
    assign mem[3068] = 12'd1027;
    assign mem[3069] = 12'd1026;
    assign mem[3070] = 12'd1025;
    assign mem[3071] = 12'd1024;
    assign mem[3072] = 12'd1023;
    assign mem[3073] = 12'd1022;
    assign mem[3074] = 12'd1021;
    assign mem[3075] = 12'd1020;
    assign mem[3076] = 12'd1019;
    assign mem[3077] = 12'd1018;
    assign mem[3078] = 12'd1017;
    assign mem[3079] = 12'd1016;
    assign mem[3080] = 12'd1015;
    assign mem[3081] = 12'd1014;
    assign mem[3082] = 12'd1013;
    assign mem[3083] = 12'd1012;
    assign mem[3084] = 12'd1011;
    assign mem[3085] = 12'd1010;
    assign mem[3086] = 12'd1009;
    assign mem[3087] = 12'd1008;
    assign mem[3088] = 12'd1007;
    assign mem[3089] = 12'd1006;
    assign mem[3090] = 12'd1005;
    assign mem[3091] = 12'd1004;
    assign mem[3092] = 12'd1003;
    assign mem[3093] = 12'd1002;
    assign mem[3094] = 12'd1001;
    assign mem[3095] = 12'd1000;
    assign mem[3096] = 12'd999;
    assign mem[3097] = 12'd998;
    assign mem[3098] = 12'd997;
    assign mem[3099] = 12'd996;
    assign mem[3100] = 12'd995;
    assign mem[3101] = 12'd994;
    assign mem[3102] = 12'd993;
    assign mem[3103] = 12'd992;
    assign mem[3104] = 12'd991;
    assign mem[3105] = 12'd990;
    assign mem[3106] = 12'd989;
    assign mem[3107] = 12'd988;
    assign mem[3108] = 12'd987;
    assign mem[3109] = 12'd986;
    assign mem[3110] = 12'd985;
    assign mem[3111] = 12'd984;
    assign mem[3112] = 12'd983;
    assign mem[3113] = 12'd982;
    assign mem[3114] = 12'd981;
    assign mem[3115] = 12'd980;
    assign mem[3116] = 12'd979;
    assign mem[3117] = 12'd978;
    assign mem[3118] = 12'd977;
    assign mem[3119] = 12'd976;
    assign mem[3120] = 12'd975;
    assign mem[3121] = 12'd974;
    assign mem[3122] = 12'd973;
    assign mem[3123] = 12'd972;
    assign mem[3124] = 12'd971;
    assign mem[3125] = 12'd970;
    assign mem[3126] = 12'd969;
    assign mem[3127] = 12'd968;
    assign mem[3128] = 12'd967;
    assign mem[3129] = 12'd966;
    assign mem[3130] = 12'd965;
    assign mem[3131] = 12'd964;
    assign mem[3132] = 12'd963;
    assign mem[3133] = 12'd962;
    assign mem[3134] = 12'd961;
    assign mem[3135] = 12'd960;
    assign mem[3136] = 12'd959;
    assign mem[3137] = 12'd958;
    assign mem[3138] = 12'd957;
    assign mem[3139] = 12'd956;
    assign mem[3140] = 12'd955;
    assign mem[3141] = 12'd954;
    assign mem[3142] = 12'd953;
    assign mem[3143] = 12'd952;
    assign mem[3144] = 12'd951;
    assign mem[3145] = 12'd950;
    assign mem[3146] = 12'd949;
    assign mem[3147] = 12'd948;
    assign mem[3148] = 12'd947;
    assign mem[3149] = 12'd946;
    assign mem[3150] = 12'd945;
    assign mem[3151] = 12'd944;
    assign mem[3152] = 12'd943;
    assign mem[3153] = 12'd942;
    assign mem[3154] = 12'd941;
    assign mem[3155] = 12'd940;
    assign mem[3156] = 12'd939;
    assign mem[3157] = 12'd938;
    assign mem[3158] = 12'd937;
    assign mem[3159] = 12'd936;
    assign mem[3160] = 12'd935;
    assign mem[3161] = 12'd934;
    assign mem[3162] = 12'd933;
    assign mem[3163] = 12'd932;
    assign mem[3164] = 12'd931;
    assign mem[3165] = 12'd930;
    assign mem[3166] = 12'd929;
    assign mem[3167] = 12'd928;
    assign mem[3168] = 12'd927;
    assign mem[3169] = 12'd926;
    assign mem[3170] = 12'd925;
    assign mem[3171] = 12'd924;
    assign mem[3172] = 12'd923;
    assign mem[3173] = 12'd922;
    assign mem[3174] = 12'd921;
    assign mem[3175] = 12'd920;
    assign mem[3176] = 12'd919;
    assign mem[3177] = 12'd918;
    assign mem[3178] = 12'd917;
    assign mem[3179] = 12'd916;
    assign mem[3180] = 12'd915;
    assign mem[3181] = 12'd914;
    assign mem[3182] = 12'd913;
    assign mem[3183] = 12'd912;
    assign mem[3184] = 12'd911;
    assign mem[3185] = 12'd910;
    assign mem[3186] = 12'd909;
    assign mem[3187] = 12'd908;
    assign mem[3188] = 12'd907;
    assign mem[3189] = 12'd906;
    assign mem[3190] = 12'd905;
    assign mem[3191] = 12'd904;
    assign mem[3192] = 12'd903;
    assign mem[3193] = 12'd902;
    assign mem[3194] = 12'd901;
    assign mem[3195] = 12'd900;
    assign mem[3196] = 12'd899;
    assign mem[3197] = 12'd898;
    assign mem[3198] = 12'd897;
    assign mem[3199] = 12'd896;
    assign mem[3200] = 12'd895;
    assign mem[3201] = 12'd894;
    assign mem[3202] = 12'd893;
    assign mem[3203] = 12'd892;
    assign mem[3204] = 12'd891;
    assign mem[3205] = 12'd890;
    assign mem[3206] = 12'd889;
    assign mem[3207] = 12'd888;
    assign mem[3208] = 12'd887;
    assign mem[3209] = 12'd886;
    assign mem[3210] = 12'd885;
    assign mem[3211] = 12'd884;
    assign mem[3212] = 12'd883;
    assign mem[3213] = 12'd882;
    assign mem[3214] = 12'd881;
    assign mem[3215] = 12'd880;
    assign mem[3216] = 12'd879;
    assign mem[3217] = 12'd878;
    assign mem[3218] = 12'd877;
    assign mem[3219] = 12'd876;
    assign mem[3220] = 12'd875;
    assign mem[3221] = 12'd874;
    assign mem[3222] = 12'd873;
    assign mem[3223] = 12'd872;
    assign mem[3224] = 12'd871;
    assign mem[3225] = 12'd870;
    assign mem[3226] = 12'd869;
    assign mem[3227] = 12'd868;
    assign mem[3228] = 12'd867;
    assign mem[3229] = 12'd866;
    assign mem[3230] = 12'd865;
    assign mem[3231] = 12'd864;
    assign mem[3232] = 12'd863;
    assign mem[3233] = 12'd862;
    assign mem[3234] = 12'd861;
    assign mem[3235] = 12'd860;
    assign mem[3236] = 12'd859;
    assign mem[3237] = 12'd858;
    assign mem[3238] = 12'd857;
    assign mem[3239] = 12'd856;
    assign mem[3240] = 12'd855;
    assign mem[3241] = 12'd854;
    assign mem[3242] = 12'd853;
    assign mem[3243] = 12'd852;
    assign mem[3244] = 12'd851;
    assign mem[3245] = 12'd850;
    assign mem[3246] = 12'd849;
    assign mem[3247] = 12'd848;
    assign mem[3248] = 12'd847;
    assign mem[3249] = 12'd846;
    assign mem[3250] = 12'd845;
    assign mem[3251] = 12'd844;
    assign mem[3252] = 12'd843;
    assign mem[3253] = 12'd842;
    assign mem[3254] = 12'd841;
    assign mem[3255] = 12'd840;
    assign mem[3256] = 12'd839;
    assign mem[3257] = 12'd838;
    assign mem[3258] = 12'd837;
    assign mem[3259] = 12'd836;
    assign mem[3260] = 12'd835;
    assign mem[3261] = 12'd834;
    assign mem[3262] = 12'd833;
    assign mem[3263] = 12'd832;
    assign mem[3264] = 12'd831;
    assign mem[3265] = 12'd830;
    assign mem[3266] = 12'd829;
    assign mem[3267] = 12'd828;
    assign mem[3268] = 12'd827;
    assign mem[3269] = 12'd826;
    assign mem[3270] = 12'd825;
    assign mem[3271] = 12'd824;
    assign mem[3272] = 12'd823;
    assign mem[3273] = 12'd822;
    assign mem[3274] = 12'd821;
    assign mem[3275] = 12'd820;
    assign mem[3276] = 12'd819;
    assign mem[3277] = 12'd818;
    assign mem[3278] = 12'd817;
    assign mem[3279] = 12'd816;
    assign mem[3280] = 12'd815;
    assign mem[3281] = 12'd814;
    assign mem[3282] = 12'd813;
    assign mem[3283] = 12'd812;
    assign mem[3284] = 12'd811;
    assign mem[3285] = 12'd810;
    assign mem[3286] = 12'd809;
    assign mem[3287] = 12'd808;
    assign mem[3288] = 12'd807;
    assign mem[3289] = 12'd806;
    assign mem[3290] = 12'd805;
    assign mem[3291] = 12'd804;
    assign mem[3292] = 12'd803;
    assign mem[3293] = 12'd802;
    assign mem[3294] = 12'd801;
    assign mem[3295] = 12'd800;
    assign mem[3296] = 12'd799;
    assign mem[3297] = 12'd798;
    assign mem[3298] = 12'd797;
    assign mem[3299] = 12'd796;
    assign mem[3300] = 12'd795;
    assign mem[3301] = 12'd794;
    assign mem[3302] = 12'd793;
    assign mem[3303] = 12'd792;
    assign mem[3304] = 12'd791;
    assign mem[3305] = 12'd790;
    assign mem[3306] = 12'd789;
    assign mem[3307] = 12'd788;
    assign mem[3308] = 12'd787;
    assign mem[3309] = 12'd786;
    assign mem[3310] = 12'd785;
    assign mem[3311] = 12'd784;
    assign mem[3312] = 12'd783;
    assign mem[3313] = 12'd782;
    assign mem[3314] = 12'd781;
    assign mem[3315] = 12'd780;
    assign mem[3316] = 12'd779;
    assign mem[3317] = 12'd778;
    assign mem[3318] = 12'd777;
    assign mem[3319] = 12'd776;
    assign mem[3320] = 12'd775;
    assign mem[3321] = 12'd774;
    assign mem[3322] = 12'd773;
    assign mem[3323] = 12'd772;
    assign mem[3324] = 12'd771;
    assign mem[3325] = 12'd770;
    assign mem[3326] = 12'd769;
    assign mem[3327] = 12'd768;
    assign mem[3328] = 12'd767;
    assign mem[3329] = 12'd766;
    assign mem[3330] = 12'd765;
    assign mem[3331] = 12'd764;
    assign mem[3332] = 12'd763;
    assign mem[3333] = 12'd762;
    assign mem[3334] = 12'd761;
    assign mem[3335] = 12'd760;
    assign mem[3336] = 12'd759;
    assign mem[3337] = 12'd758;
    assign mem[3338] = 12'd757;
    assign mem[3339] = 12'd756;
    assign mem[3340] = 12'd755;
    assign mem[3341] = 12'd754;
    assign mem[3342] = 12'd753;
    assign mem[3343] = 12'd752;
    assign mem[3344] = 12'd751;
    assign mem[3345] = 12'd750;
    assign mem[3346] = 12'd749;
    assign mem[3347] = 12'd748;
    assign mem[3348] = 12'd747;
    assign mem[3349] = 12'd746;
    assign mem[3350] = 12'd745;
    assign mem[3351] = 12'd744;
    assign mem[3352] = 12'd743;
    assign mem[3353] = 12'd742;
    assign mem[3354] = 12'd741;
    assign mem[3355] = 12'd740;
    assign mem[3356] = 12'd739;
    assign mem[3357] = 12'd738;
    assign mem[3358] = 12'd737;
    assign mem[3359] = 12'd736;
    assign mem[3360] = 12'd735;
    assign mem[3361] = 12'd734;
    assign mem[3362] = 12'd733;
    assign mem[3363] = 12'd732;
    assign mem[3364] = 12'd731;
    assign mem[3365] = 12'd730;
    assign mem[3366] = 12'd729;
    assign mem[3367] = 12'd728;
    assign mem[3368] = 12'd727;
    assign mem[3369] = 12'd726;
    assign mem[3370] = 12'd725;
    assign mem[3371] = 12'd724;
    assign mem[3372] = 12'd723;
    assign mem[3373] = 12'd722;
    assign mem[3374] = 12'd721;
    assign mem[3375] = 12'd720;
    assign mem[3376] = 12'd719;
    assign mem[3377] = 12'd718;
    assign mem[3378] = 12'd717;
    assign mem[3379] = 12'd716;
    assign mem[3380] = 12'd715;
    assign mem[3381] = 12'd714;
    assign mem[3382] = 12'd713;
    assign mem[3383] = 12'd712;
    assign mem[3384] = 12'd711;
    assign mem[3385] = 12'd710;
    assign mem[3386] = 12'd709;
    assign mem[3387] = 12'd708;
    assign mem[3388] = 12'd707;
    assign mem[3389] = 12'd706;
    assign mem[3390] = 12'd705;
    assign mem[3391] = 12'd704;
    assign mem[3392] = 12'd703;
    assign mem[3393] = 12'd702;
    assign mem[3394] = 12'd701;
    assign mem[3395] = 12'd700;
    assign mem[3396] = 12'd699;
    assign mem[3397] = 12'd698;
    assign mem[3398] = 12'd697;
    assign mem[3399] = 12'd696;
    assign mem[3400] = 12'd695;
    assign mem[3401] = 12'd694;
    assign mem[3402] = 12'd693;
    assign mem[3403] = 12'd692;
    assign mem[3404] = 12'd691;
    assign mem[3405] = 12'd690;
    assign mem[3406] = 12'd689;
    assign mem[3407] = 12'd688;
    assign mem[3408] = 12'd687;
    assign mem[3409] = 12'd686;
    assign mem[3410] = 12'd685;
    assign mem[3411] = 12'd684;
    assign mem[3412] = 12'd683;
    assign mem[3413] = 12'd682;
    assign mem[3414] = 12'd681;
    assign mem[3415] = 12'd680;
    assign mem[3416] = 12'd679;
    assign mem[3417] = 12'd678;
    assign mem[3418] = 12'd677;
    assign mem[3419] = 12'd676;
    assign mem[3420] = 12'd675;
    assign mem[3421] = 12'd674;
    assign mem[3422] = 12'd673;
    assign mem[3423] = 12'd672;
    assign mem[3424] = 12'd671;
    assign mem[3425] = 12'd670;
    assign mem[3426] = 12'd669;
    assign mem[3427] = 12'd668;
    assign mem[3428] = 12'd667;
    assign mem[3429] = 12'd666;
    assign mem[3430] = 12'd665;
    assign mem[3431] = 12'd664;
    assign mem[3432] = 12'd663;
    assign mem[3433] = 12'd662;
    assign mem[3434] = 12'd661;
    assign mem[3435] = 12'd660;
    assign mem[3436] = 12'd659;
    assign mem[3437] = 12'd658;
    assign mem[3438] = 12'd657;
    assign mem[3439] = 12'd656;
    assign mem[3440] = 12'd655;
    assign mem[3441] = 12'd654;
    assign mem[3442] = 12'd653;
    assign mem[3443] = 12'd652;
    assign mem[3444] = 12'd651;
    assign mem[3445] = 12'd650;
    assign mem[3446] = 12'd649;
    assign mem[3447] = 12'd648;
    assign mem[3448] = 12'd647;
    assign mem[3449] = 12'd646;
    assign mem[3450] = 12'd645;
    assign mem[3451] = 12'd644;
    assign mem[3452] = 12'd643;
    assign mem[3453] = 12'd642;
    assign mem[3454] = 12'd641;
    assign mem[3455] = 12'd640;
    assign mem[3456] = 12'd639;
    assign mem[3457] = 12'd638;
    assign mem[3458] = 12'd637;
    assign mem[3459] = 12'd636;
    assign mem[3460] = 12'd635;
    assign mem[3461] = 12'd634;
    assign mem[3462] = 12'd633;
    assign mem[3463] = 12'd632;
    assign mem[3464] = 12'd631;
    assign mem[3465] = 12'd630;
    assign mem[3466] = 12'd629;
    assign mem[3467] = 12'd628;
    assign mem[3468] = 12'd627;
    assign mem[3469] = 12'd626;
    assign mem[3470] = 12'd625;
    assign mem[3471] = 12'd624;
    assign mem[3472] = 12'd623;
    assign mem[3473] = 12'd622;
    assign mem[3474] = 12'd621;
    assign mem[3475] = 12'd620;
    assign mem[3476] = 12'd619;
    assign mem[3477] = 12'd618;
    assign mem[3478] = 12'd617;
    assign mem[3479] = 12'd616;
    assign mem[3480] = 12'd615;
    assign mem[3481] = 12'd614;
    assign mem[3482] = 12'd613;
    assign mem[3483] = 12'd612;
    assign mem[3484] = 12'd611;
    assign mem[3485] = 12'd610;
    assign mem[3486] = 12'd609;
    assign mem[3487] = 12'd608;
    assign mem[3488] = 12'd607;
    assign mem[3489] = 12'd606;
    assign mem[3490] = 12'd605;
    assign mem[3491] = 12'd604;
    assign mem[3492] = 12'd603;
    assign mem[3493] = 12'd602;
    assign mem[3494] = 12'd601;
    assign mem[3495] = 12'd600;
    assign mem[3496] = 12'd599;
    assign mem[3497] = 12'd598;
    assign mem[3498] = 12'd597;
    assign mem[3499] = 12'd596;
    assign mem[3500] = 12'd595;
    assign mem[3501] = 12'd594;
    assign mem[3502] = 12'd593;
    assign mem[3503] = 12'd592;
    assign mem[3504] = 12'd591;
    assign mem[3505] = 12'd590;
    assign mem[3506] = 12'd589;
    assign mem[3507] = 12'd588;
    assign mem[3508] = 12'd587;
    assign mem[3509] = 12'd586;
    assign mem[3510] = 12'd585;
    assign mem[3511] = 12'd584;
    assign mem[3512] = 12'd583;
    assign mem[3513] = 12'd582;
    assign mem[3514] = 12'd581;
    assign mem[3515] = 12'd580;
    assign mem[3516] = 12'd579;
    assign mem[3517] = 12'd578;
    assign mem[3518] = 12'd577;
    assign mem[3519] = 12'd576;
    assign mem[3520] = 12'd575;
    assign mem[3521] = 12'd574;
    assign mem[3522] = 12'd573;
    assign mem[3523] = 12'd572;
    assign mem[3524] = 12'd571;
    assign mem[3525] = 12'd570;
    assign mem[3526] = 12'd569;
    assign mem[3527] = 12'd568;
    assign mem[3528] = 12'd567;
    assign mem[3529] = 12'd566;
    assign mem[3530] = 12'd565;
    assign mem[3531] = 12'd564;
    assign mem[3532] = 12'd563;
    assign mem[3533] = 12'd562;
    assign mem[3534] = 12'd561;
    assign mem[3535] = 12'd560;
    assign mem[3536] = 12'd559;
    assign mem[3537] = 12'd558;
    assign mem[3538] = 12'd557;
    assign mem[3539] = 12'd556;
    assign mem[3540] = 12'd555;
    assign mem[3541] = 12'd554;
    assign mem[3542] = 12'd553;
    assign mem[3543] = 12'd552;
    assign mem[3544] = 12'd551;
    assign mem[3545] = 12'd550;
    assign mem[3546] = 12'd549;
    assign mem[3547] = 12'd548;
    assign mem[3548] = 12'd547;
    assign mem[3549] = 12'd546;
    assign mem[3550] = 12'd545;
    assign mem[3551] = 12'd544;
    assign mem[3552] = 12'd543;
    assign mem[3553] = 12'd542;
    assign mem[3554] = 12'd541;
    assign mem[3555] = 12'd540;
    assign mem[3556] = 12'd539;
    assign mem[3557] = 12'd538;
    assign mem[3558] = 12'd537;
    assign mem[3559] = 12'd536;
    assign mem[3560] = 12'd535;
    assign mem[3561] = 12'd534;
    assign mem[3562] = 12'd533;
    assign mem[3563] = 12'd532;
    assign mem[3564] = 12'd531;
    assign mem[3565] = 12'd530;
    assign mem[3566] = 12'd529;
    assign mem[3567] = 12'd528;
    assign mem[3568] = 12'd527;
    assign mem[3569] = 12'd526;
    assign mem[3570] = 12'd525;
    assign mem[3571] = 12'd524;
    assign mem[3572] = 12'd523;
    assign mem[3573] = 12'd522;
    assign mem[3574] = 12'd521;
    assign mem[3575] = 12'd520;
    assign mem[3576] = 12'd519;
    assign mem[3577] = 12'd518;
    assign mem[3578] = 12'd517;
    assign mem[3579] = 12'd516;
    assign mem[3580] = 12'd515;
    assign mem[3581] = 12'd514;
    assign mem[3582] = 12'd513;
    assign mem[3583] = 12'd512;
    assign mem[3584] = 12'd511;
    assign mem[3585] = 12'd510;
    assign mem[3586] = 12'd509;
    assign mem[3587] = 12'd508;
    assign mem[3588] = 12'd507;
    assign mem[3589] = 12'd506;
    assign mem[3590] = 12'd505;
    assign mem[3591] = 12'd504;
    assign mem[3592] = 12'd503;
    assign mem[3593] = 12'd502;
    assign mem[3594] = 12'd501;
    assign mem[3595] = 12'd500;
    assign mem[3596] = 12'd499;
    assign mem[3597] = 12'd498;
    assign mem[3598] = 12'd497;
    assign mem[3599] = 12'd496;
    assign mem[3600] = 12'd495;
    assign mem[3601] = 12'd494;
    assign mem[3602] = 12'd493;
    assign mem[3603] = 12'd492;
    assign mem[3604] = 12'd491;
    assign mem[3605] = 12'd490;
    assign mem[3606] = 12'd489;
    assign mem[3607] = 12'd488;
    assign mem[3608] = 12'd487;
    assign mem[3609] = 12'd486;
    assign mem[3610] = 12'd485;
    assign mem[3611] = 12'd484;
    assign mem[3612] = 12'd483;
    assign mem[3613] = 12'd482;
    assign mem[3614] = 12'd481;
    assign mem[3615] = 12'd480;
    assign mem[3616] = 12'd479;
    assign mem[3617] = 12'd478;
    assign mem[3618] = 12'd477;
    assign mem[3619] = 12'd476;
    assign mem[3620] = 12'd475;
    assign mem[3621] = 12'd474;
    assign mem[3622] = 12'd473;
    assign mem[3623] = 12'd472;
    assign mem[3624] = 12'd471;
    assign mem[3625] = 12'd470;
    assign mem[3626] = 12'd469;
    assign mem[3627] = 12'd468;
    assign mem[3628] = 12'd467;
    assign mem[3629] = 12'd466;
    assign mem[3630] = 12'd465;
    assign mem[3631] = 12'd464;
    assign mem[3632] = 12'd463;
    assign mem[3633] = 12'd462;
    assign mem[3634] = 12'd461;
    assign mem[3635] = 12'd460;
    assign mem[3636] = 12'd459;
    assign mem[3637] = 12'd458;
    assign mem[3638] = 12'd457;
    assign mem[3639] = 12'd456;
    assign mem[3640] = 12'd455;
    assign mem[3641] = 12'd454;
    assign mem[3642] = 12'd453;
    assign mem[3643] = 12'd452;
    assign mem[3644] = 12'd451;
    assign mem[3645] = 12'd450;
    assign mem[3646] = 12'd449;
    assign mem[3647] = 12'd448;
    assign mem[3648] = 12'd447;
    assign mem[3649] = 12'd446;
    assign mem[3650] = 12'd445;
    assign mem[3651] = 12'd444;
    assign mem[3652] = 12'd443;
    assign mem[3653] = 12'd442;
    assign mem[3654] = 12'd441;
    assign mem[3655] = 12'd440;
    assign mem[3656] = 12'd439;
    assign mem[3657] = 12'd438;
    assign mem[3658] = 12'd437;
    assign mem[3659] = 12'd436;
    assign mem[3660] = 12'd435;
    assign mem[3661] = 12'd434;
    assign mem[3662] = 12'd433;
    assign mem[3663] = 12'd432;
    assign mem[3664] = 12'd431;
    assign mem[3665] = 12'd430;
    assign mem[3666] = 12'd429;
    assign mem[3667] = 12'd428;
    assign mem[3668] = 12'd427;
    assign mem[3669] = 12'd426;
    assign mem[3670] = 12'd425;
    assign mem[3671] = 12'd424;
    assign mem[3672] = 12'd423;
    assign mem[3673] = 12'd422;
    assign mem[3674] = 12'd421;
    assign mem[3675] = 12'd420;
    assign mem[3676] = 12'd419;
    assign mem[3677] = 12'd418;
    assign mem[3678] = 12'd417;
    assign mem[3679] = 12'd416;
    assign mem[3680] = 12'd415;
    assign mem[3681] = 12'd414;
    assign mem[3682] = 12'd413;
    assign mem[3683] = 12'd412;
    assign mem[3684] = 12'd411;
    assign mem[3685] = 12'd410;
    assign mem[3686] = 12'd409;
    assign mem[3687] = 12'd408;
    assign mem[3688] = 12'd407;
    assign mem[3689] = 12'd406;
    assign mem[3690] = 12'd405;
    assign mem[3691] = 12'd404;
    assign mem[3692] = 12'd403;
    assign mem[3693] = 12'd402;
    assign mem[3694] = 12'd401;
    assign mem[3695] = 12'd400;
    assign mem[3696] = 12'd399;
    assign mem[3697] = 12'd398;
    assign mem[3698] = 12'd397;
    assign mem[3699] = 12'd396;
    assign mem[3700] = 12'd395;
    assign mem[3701] = 12'd394;
    assign mem[3702] = 12'd393;
    assign mem[3703] = 12'd392;
    assign mem[3704] = 12'd391;
    assign mem[3705] = 12'd390;
    assign mem[3706] = 12'd389;
    assign mem[3707] = 12'd388;
    assign mem[3708] = 12'd387;
    assign mem[3709] = 12'd386;
    assign mem[3710] = 12'd385;
    assign mem[3711] = 12'd384;
    assign mem[3712] = 12'd383;
    assign mem[3713] = 12'd382;
    assign mem[3714] = 12'd381;
    assign mem[3715] = 12'd380;
    assign mem[3716] = 12'd379;
    assign mem[3717] = 12'd378;
    assign mem[3718] = 12'd377;
    assign mem[3719] = 12'd376;
    assign mem[3720] = 12'd375;
    assign mem[3721] = 12'd374;
    assign mem[3722] = 12'd373;
    assign mem[3723] = 12'd372;
    assign mem[3724] = 12'd371;
    assign mem[3725] = 12'd370;
    assign mem[3726] = 12'd369;
    assign mem[3727] = 12'd368;
    assign mem[3728] = 12'd367;
    assign mem[3729] = 12'd366;
    assign mem[3730] = 12'd365;
    assign mem[3731] = 12'd364;
    assign mem[3732] = 12'd363;
    assign mem[3733] = 12'd362;
    assign mem[3734] = 12'd361;
    assign mem[3735] = 12'd360;
    assign mem[3736] = 12'd359;
    assign mem[3737] = 12'd358;
    assign mem[3738] = 12'd357;
    assign mem[3739] = 12'd356;
    assign mem[3740] = 12'd355;
    assign mem[3741] = 12'd354;
    assign mem[3742] = 12'd353;
    assign mem[3743] = 12'd352;
    assign mem[3744] = 12'd351;
    assign mem[3745] = 12'd350;
    assign mem[3746] = 12'd349;
    assign mem[3747] = 12'd348;
    assign mem[3748] = 12'd347;
    assign mem[3749] = 12'd346;
    assign mem[3750] = 12'd345;
    assign mem[3751] = 12'd344;
    assign mem[3752] = 12'd343;
    assign mem[3753] = 12'd342;
    assign mem[3754] = 12'd341;
    assign mem[3755] = 12'd340;
    assign mem[3756] = 12'd339;
    assign mem[3757] = 12'd338;
    assign mem[3758] = 12'd337;
    assign mem[3759] = 12'd336;
    assign mem[3760] = 12'd335;
    assign mem[3761] = 12'd334;
    assign mem[3762] = 12'd333;
    assign mem[3763] = 12'd332;
    assign mem[3764] = 12'd331;
    assign mem[3765] = 12'd330;
    assign mem[3766] = 12'd329;
    assign mem[3767] = 12'd328;
    assign mem[3768] = 12'd327;
    assign mem[3769] = 12'd326;
    assign mem[3770] = 12'd325;
    assign mem[3771] = 12'd324;
    assign mem[3772] = 12'd323;
    assign mem[3773] = 12'd322;
    assign mem[3774] = 12'd321;
    assign mem[3775] = 12'd320;
    assign mem[3776] = 12'd319;
    assign mem[3777] = 12'd318;
    assign mem[3778] = 12'd317;
    assign mem[3779] = 12'd316;
    assign mem[3780] = 12'd315;
    assign mem[3781] = 12'd314;
    assign mem[3782] = 12'd313;
    assign mem[3783] = 12'd312;
    assign mem[3784] = 12'd311;
    assign mem[3785] = 12'd310;
    assign mem[3786] = 12'd309;
    assign mem[3787] = 12'd308;
    assign mem[3788] = 12'd307;
    assign mem[3789] = 12'd306;
    assign mem[3790] = 12'd305;
    assign mem[3791] = 12'd304;
    assign mem[3792] = 12'd303;
    assign mem[3793] = 12'd302;
    assign mem[3794] = 12'd301;
    assign mem[3795] = 12'd300;
    assign mem[3796] = 12'd299;
    assign mem[3797] = 12'd298;
    assign mem[3798] = 12'd297;
    assign mem[3799] = 12'd296;
    assign mem[3800] = 12'd295;
    assign mem[3801] = 12'd294;
    assign mem[3802] = 12'd293;
    assign mem[3803] = 12'd292;
    assign mem[3804] = 12'd291;
    assign mem[3805] = 12'd290;
    assign mem[3806] = 12'd289;
    assign mem[3807] = 12'd288;
    assign mem[3808] = 12'd287;
    assign mem[3809] = 12'd286;
    assign mem[3810] = 12'd285;
    assign mem[3811] = 12'd284;
    assign mem[3812] = 12'd283;
    assign mem[3813] = 12'd282;
    assign mem[3814] = 12'd281;
    assign mem[3815] = 12'd280;
    assign mem[3816] = 12'd279;
    assign mem[3817] = 12'd278;
    assign mem[3818] = 12'd277;
    assign mem[3819] = 12'd276;
    assign mem[3820] = 12'd275;
    assign mem[3821] = 12'd274;
    assign mem[3822] = 12'd273;
    assign mem[3823] = 12'd272;
    assign mem[3824] = 12'd271;
    assign mem[3825] = 12'd270;
    assign mem[3826] = 12'd269;
    assign mem[3827] = 12'd268;
    assign mem[3828] = 12'd267;
    assign mem[3829] = 12'd266;
    assign mem[3830] = 12'd265;
    assign mem[3831] = 12'd264;
    assign mem[3832] = 12'd263;
    assign mem[3833] = 12'd262;
    assign mem[3834] = 12'd261;
    assign mem[3835] = 12'd260;
    assign mem[3836] = 12'd259;
    assign mem[3837] = 12'd258;
    assign mem[3838] = 12'd257;
    assign mem[3839] = 12'd256;
    assign mem[3840] = 12'd255;
    assign mem[3841] = 12'd254;
    assign mem[3842] = 12'd253;
    assign mem[3843] = 12'd252;
    assign mem[3844] = 12'd251;
    assign mem[3845] = 12'd250;
    assign mem[3846] = 12'd249;
    assign mem[3847] = 12'd248;
    assign mem[3848] = 12'd247;
    assign mem[3849] = 12'd246;
    assign mem[3850] = 12'd245;
    assign mem[3851] = 12'd244;
    assign mem[3852] = 12'd243;
    assign mem[3853] = 12'd242;
    assign mem[3854] = 12'd241;
    assign mem[3855] = 12'd240;
    assign mem[3856] = 12'd239;
    assign mem[3857] = 12'd238;
    assign mem[3858] = 12'd237;
    assign mem[3859] = 12'd236;
    assign mem[3860] = 12'd235;
    assign mem[3861] = 12'd234;
    assign mem[3862] = 12'd233;
    assign mem[3863] = 12'd232;
    assign mem[3864] = 12'd231;
    assign mem[3865] = 12'd230;
    assign mem[3866] = 12'd229;
    assign mem[3867] = 12'd228;
    assign mem[3868] = 12'd227;
    assign mem[3869] = 12'd226;
    assign mem[3870] = 12'd225;
    assign mem[3871] = 12'd224;
    assign mem[3872] = 12'd223;
    assign mem[3873] = 12'd222;
    assign mem[3874] = 12'd221;
    assign mem[3875] = 12'd220;
    assign mem[3876] = 12'd219;
    assign mem[3877] = 12'd218;
    assign mem[3878] = 12'd217;
    assign mem[3879] = 12'd216;
    assign mem[3880] = 12'd215;
    assign mem[3881] = 12'd214;
    assign mem[3882] = 12'd213;
    assign mem[3883] = 12'd212;
    assign mem[3884] = 12'd211;
    assign mem[3885] = 12'd210;
    assign mem[3886] = 12'd209;
    assign mem[3887] = 12'd208;
    assign mem[3888] = 12'd207;
    assign mem[3889] = 12'd206;
    assign mem[3890] = 12'd205;
    assign mem[3891] = 12'd204;
    assign mem[3892] = 12'd203;
    assign mem[3893] = 12'd202;
    assign mem[3894] = 12'd201;
    assign mem[3895] = 12'd200;
    assign mem[3896] = 12'd199;
    assign mem[3897] = 12'd198;
    assign mem[3898] = 12'd197;
    assign mem[3899] = 12'd196;
    assign mem[3900] = 12'd195;
    assign mem[3901] = 12'd194;
    assign mem[3902] = 12'd193;
    assign mem[3903] = 12'd192;
    assign mem[3904] = 12'd191;
    assign mem[3905] = 12'd190;
    assign mem[3906] = 12'd189;
    assign mem[3907] = 12'd188;
    assign mem[3908] = 12'd187;
    assign mem[3909] = 12'd186;
    assign mem[3910] = 12'd185;
    assign mem[3911] = 12'd184;
    assign mem[3912] = 12'd183;
    assign mem[3913] = 12'd182;
    assign mem[3914] = 12'd181;
    assign mem[3915] = 12'd180;
    assign mem[3916] = 12'd179;
    assign mem[3917] = 12'd178;
    assign mem[3918] = 12'd177;
    assign mem[3919] = 12'd176;
    assign mem[3920] = 12'd175;
    assign mem[3921] = 12'd174;
    assign mem[3922] = 12'd173;
    assign mem[3923] = 12'd172;
    assign mem[3924] = 12'd171;
    assign mem[3925] = 12'd170;
    assign mem[3926] = 12'd169;
    assign mem[3927] = 12'd168;
    assign mem[3928] = 12'd167;
    assign mem[3929] = 12'd166;
    assign mem[3930] = 12'd165;
    assign mem[3931] = 12'd164;
    assign mem[3932] = 12'd163;
    assign mem[3933] = 12'd162;
    assign mem[3934] = 12'd161;
    assign mem[3935] = 12'd160;
    assign mem[3936] = 12'd159;
    assign mem[3937] = 12'd158;
    assign mem[3938] = 12'd157;
    assign mem[3939] = 12'd156;
    assign mem[3940] = 12'd155;
    assign mem[3941] = 12'd154;
    assign mem[3942] = 12'd153;
    assign mem[3943] = 12'd152;
    assign mem[3944] = 12'd151;
    assign mem[3945] = 12'd150;
    assign mem[3946] = 12'd149;
    assign mem[3947] = 12'd148;
    assign mem[3948] = 12'd147;
    assign mem[3949] = 12'd146;
    assign mem[3950] = 12'd145;
    assign mem[3951] = 12'd144;
    assign mem[3952] = 12'd143;
    assign mem[3953] = 12'd142;
    assign mem[3954] = 12'd141;
    assign mem[3955] = 12'd140;
    assign mem[3956] = 12'd139;
    assign mem[3957] = 12'd138;
    assign mem[3958] = 12'd137;
    assign mem[3959] = 12'd136;
    assign mem[3960] = 12'd135;
    assign mem[3961] = 12'd134;
    assign mem[3962] = 12'd133;
    assign mem[3963] = 12'd132;
    assign mem[3964] = 12'd131;
    assign mem[3965] = 12'd130;
    assign mem[3966] = 12'd129;
    assign mem[3967] = 12'd128;
    assign mem[3968] = 12'd127;
    assign mem[3969] = 12'd126;
    assign mem[3970] = 12'd125;
    assign mem[3971] = 12'd124;
    assign mem[3972] = 12'd123;
    assign mem[3973] = 12'd122;
    assign mem[3974] = 12'd121;
    assign mem[3975] = 12'd120;
    assign mem[3976] = 12'd119;
    assign mem[3977] = 12'd118;
    assign mem[3978] = 12'd117;
    assign mem[3979] = 12'd116;
    assign mem[3980] = 12'd115;
    assign mem[3981] = 12'd114;
    assign mem[3982] = 12'd113;
    assign mem[3983] = 12'd112;
    assign mem[3984] = 12'd111;
    assign mem[3985] = 12'd110;
    assign mem[3986] = 12'd109;
    assign mem[3987] = 12'd108;
    assign mem[3988] = 12'd107;
    assign mem[3989] = 12'd106;
    assign mem[3990] = 12'd105;
    assign mem[3991] = 12'd104;
    assign mem[3992] = 12'd103;
    assign mem[3993] = 12'd102;
    assign mem[3994] = 12'd101;
    assign mem[3995] = 12'd100;
    assign mem[3996] = 12'd99;
    assign mem[3997] = 12'd98;
    assign mem[3998] = 12'd97;
    assign mem[3999] = 12'd96;
    assign mem[4000] = 12'd95;
    assign mem[4001] = 12'd94;
    assign mem[4002] = 12'd93;
    assign mem[4003] = 12'd92;
    assign mem[4004] = 12'd91;
    assign mem[4005] = 12'd90;
    assign mem[4006] = 12'd89;
    assign mem[4007] = 12'd88;
    assign mem[4008] = 12'd87;
    assign mem[4009] = 12'd86;
    assign mem[4010] = 12'd85;
    assign mem[4011] = 12'd84;
    assign mem[4012] = 12'd83;
    assign mem[4013] = 12'd82;
    assign mem[4014] = 12'd81;
    assign mem[4015] = 12'd80;
    assign mem[4016] = 12'd79;
    assign mem[4017] = 12'd78;
    assign mem[4018] = 12'd77;
    assign mem[4019] = 12'd76;
    assign mem[4020] = 12'd75;
    assign mem[4021] = 12'd74;
    assign mem[4022] = 12'd73;
    assign mem[4023] = 12'd72;
    assign mem[4024] = 12'd71;
    assign mem[4025] = 12'd70;
    assign mem[4026] = 12'd69;
    assign mem[4027] = 12'd68;
    assign mem[4028] = 12'd67;
    assign mem[4029] = 12'd66;
    assign mem[4030] = 12'd65;
    assign mem[4031] = 12'd64;
    assign mem[4032] = 12'd63;
    assign mem[4033] = 12'd62;
    assign mem[4034] = 12'd61;
    assign mem[4035] = 12'd60;
    assign mem[4036] = 12'd59;
    assign mem[4037] = 12'd58;
    assign mem[4038] = 12'd57;
    assign mem[4039] = 12'd56;
    assign mem[4040] = 12'd55;
    assign mem[4041] = 12'd54;
    assign mem[4042] = 12'd53;
    assign mem[4043] = 12'd52;
    assign mem[4044] = 12'd51;
    assign mem[4045] = 12'd50;
    assign mem[4046] = 12'd49;
    assign mem[4047] = 12'd48;
    assign mem[4048] = 12'd47;
    assign mem[4049] = 12'd46;
    assign mem[4050] = 12'd45;
    assign mem[4051] = 12'd44;
    assign mem[4052] = 12'd43;
    assign mem[4053] = 12'd42;
    assign mem[4054] = 12'd41;
    assign mem[4055] = 12'd40;
    assign mem[4056] = 12'd39;
    assign mem[4057] = 12'd38;
    assign mem[4058] = 12'd37;
    assign mem[4059] = 12'd36;
    assign mem[4060] = 12'd35;
    assign mem[4061] = 12'd34;
    assign mem[4062] = 12'd33;
    assign mem[4063] = 12'd32;
    assign mem[4064] = 12'd31;
    assign mem[4065] = 12'd30;
    assign mem[4066] = 12'd29;
    assign mem[4067] = 12'd28;
    assign mem[4068] = 12'd27;
    assign mem[4069] = 12'd26;
    assign mem[4070] = 12'd25;
    assign mem[4071] = 12'd24;
    assign mem[4072] = 12'd23;
    assign mem[4073] = 12'd22;
    assign mem[4074] = 12'd21;
    assign mem[4075] = 12'd20;
    assign mem[4076] = 12'd19;
    assign mem[4077] = 12'd18;
    assign mem[4078] = 12'd17;
    assign mem[4079] = 12'd16;
    assign mem[4080] = 12'd15;
    assign mem[4081] = 12'd14;
    assign mem[4082] = 12'd13;
    assign mem[4083] = 12'd12;
    assign mem[4084] = 12'd11;
    assign mem[4085] = 12'd10;
    assign mem[4086] = 12'd9;
    assign mem[4087] = 12'd8;
    assign mem[4088] = 12'd7;
    assign mem[4089] = 12'd6;
    assign mem[4090] = 12'd5;
    assign mem[4091] = 12'd4;
    assign mem[4092] = 12'd3;
    assign mem[4093] = 12'd2;
    assign mem[4094] = 12'd1;
    assign mem[4095] = 12'd0;


endmodule